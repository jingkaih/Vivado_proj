module ALU(
  input         clock,
  input         reset,
  input  [8:0]  io_opcode,
  input  [63:0] io_in_a,
  input  [63:0] io_in_b,
  output [63:0] io_out_a,
  output [63:0] io_out_b,
  input         io_validin_a,
  output        io_validout_a
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] snapshot_a; // @[ALU.scala 25:27]
  reg [63:0] snapshot_b; // @[ALU.scala 26:27]
  reg  snapshot_valid_a; // @[ALU.scala 28:33]
  reg [63:0] temp_result_a; // @[ALU.scala 33:30]
  reg [63:0] temp_result_b; // @[ALU.scala 34:30]
  reg  temp_valid_a; // @[ALU.scala 37:29]
  wire  opcode_0 = io_opcode[0]; // @[ALU.scala 41:34]
  wire  opcode_1 = io_opcode[1]; // @[ALU.scala 41:34]
  wire  opcode_2 = io_opcode[2]; // @[ALU.scala 41:34]
  wire  opcode_3 = io_opcode[3]; // @[ALU.scala 41:34]
  wire  opcode_4 = io_opcode[4]; // @[ALU.scala 41:34]
  wire  opcode_5 = io_opcode[5]; // @[ALU.scala 41:34]
  wire  opcode_6 = io_opcode[6]; // @[ALU.scala 41:34]
  wire  opcode_7 = io_opcode[7]; // @[ALU.scala 41:34]
  wire  opcode_8 = io_opcode[8]; // @[ALU.scala 41:34]
  wire  _T_1 = ~opcode_7; // @[ALU.scala 51:39]
  wire  _T_5 = opcode_6 & opcode_5; // @[ALU.scala 52:28]
  wire  _T_26 = ~opcode_4; // @[ALU.scala 93:20]
  wire  _T_27 = ~opcode_3; // @[ALU.scala 93:41]
  wire  _T_28 = ~opcode_4 & ~opcode_3; // @[ALU.scala 93:28]
  wire [63:0] _gate_a_T = ~io_in_a; // @[ALU.scala 94:17]
  wire  _T_31 = opcode_4 & _T_27; // @[ALU.scala 98:34]
  wire [63:0] _gate_a_T_1 = ~snapshot_a; // @[ALU.scala 99:17]
  wire  _T_34 = _T_26 & opcode_3; // @[ALU.scala 103:34]
  wire [63:0] _GEN_18 = _T_26 & opcode_3 ? _gate_a_T : _gate_a_T_1; // @[ALU.scala 103:55 ALU.scala 104:14 ALU.scala 109:14]
  wire [63:0] _GEN_22 = opcode_4 & _T_27 ? _gate_a_T_1 : _GEN_18; // @[ALU.scala 98:55 ALU.scala 99:14]
  wire [63:0] _GEN_26 = ~opcode_4 & ~opcode_3 ? _gate_a_T : _GEN_22; // @[ALU.scala 93:49 ALU.scala 94:14]
  wire  _T_38 = ~opcode_5; // @[ALU.scala 114:66]
  wire [63:0] _GEN_30 = _T_34 ? io_in_a : snapshot_a; // @[ALU.scala 125:55 ALU.scala 126:14 ALU.scala 131:14]
  wire [63:0] _GEN_34 = _T_31 ? snapshot_a : _GEN_30; // @[ALU.scala 120:55 ALU.scala 121:14]
  wire [63:0] _GEN_38 = _T_28 ? io_in_a : _GEN_34; // @[ALU.scala 115:49 ALU.scala 116:14]
  wire [63:0] _GEN_54 = opcode_8 & opcode_6 & ~opcode_5 ? _GEN_38 : _GEN_38; // @[ALU.scala 114:74]
  wire [63:0] gate_a = opcode_8 & ~opcode_6 & opcode_5 ? _GEN_26 : _GEN_54; // @[ALU.scala 92:68]
  wire [63:0] _GEN_23 = opcode_4 & _T_27 ? io_in_b : snapshot_b; // @[ALU.scala 98:55 ALU.scala 100:14]
  wire [63:0] _GEN_27 = ~opcode_4 & ~opcode_3 ? io_in_b : _GEN_23; // @[ALU.scala 93:49 ALU.scala 95:14]
  wire [63:0] _gate_b_T = ~io_in_b; // @[ALU.scala 117:17]
  wire [63:0] _gate_b_T_2 = ~snapshot_b; // @[ALU.scala 127:17]
  wire [63:0] _GEN_31 = _T_34 ? _gate_b_T_2 : _gate_b_T_2; // @[ALU.scala 125:55 ALU.scala 127:14 ALU.scala 132:14]
  wire [63:0] _GEN_35 = _T_31 ? _gate_b_T : _GEN_31; // @[ALU.scala 120:55 ALU.scala 122:14]
  wire [63:0] _GEN_39 = _T_28 ? _gate_b_T : _GEN_35; // @[ALU.scala 115:49 ALU.scala 117:14]
  wire [63:0] _GEN_55 = opcode_8 & opcode_6 & ~opcode_5 ? _GEN_39 : _GEN_27; // @[ALU.scala 114:74]
  wire [63:0] gate_b = opcode_8 & ~opcode_6 & opcode_5 ? _GEN_27 : _GEN_55; // @[ALU.scala 92:68]
  wire [63:0] _temp_result_a_T = gate_a & gate_b; // @[ALU.scala 53:33]
  wire [63:0] _temp_result_a_T_1 = ~_temp_result_a_T; // @[ALU.scala 53:24]
  wire [63:0] _temp_result_a_T_3 = gate_a | gate_b; // @[ALU.scala 61:33]
  wire [63:0] _temp_result_a_T_4 = ~_temp_result_a_T_3; // @[ALU.scala 61:24]
  wire  _T_12 = ~opcode_8; // @[ALU.scala 67:24]
  wire [63:0] _temp_result_a_T_6 = gate_a ^ gate_b; // @[ALU.scala 69:33]
  wire [63:0] _temp_result_a_T_7 = ~_temp_result_a_T_6; // @[ALU.scala 69:24]
  wire [63:0] _GEN_4 = opcode_5 ? _temp_result_a_T_7 : _temp_result_a_T_6; // @[ALU.scala 68:28 ALU.scala 69:21 ALU.scala 72:21]
  wire  _T_18 = _T_12 & _T_1; // @[ALU.scala 75:32]
  wire [63:0] _temp_result_a_T_9 = ~gate_a; // @[ALU.scala 80:24]
  wire [63:0] _GEN_6 = opcode_5 ? _temp_result_a_T_9 : temp_result_a; // @[ALU.scala 79:34 ALU.scala 80:21 ALU.scala 33:30]
  wire [63:0] _GEN_7 = opcode_5 ? gate_b : temp_result_b; // @[ALU.scala 79:34 ALU.scala 81:21 ALU.scala 34:30]
  wire [63:0] _GEN_8 = _T_38 ? gate_a : _GEN_6; // @[ALU.scala 76:28 ALU.scala 77:21]
  wire [63:0] _GEN_9 = _T_38 ? gate_b : _GEN_7; // @[ALU.scala 76:28 ALU.scala 78:21]
  wire [63:0] _GEN_10 = _T_12 & _T_1 ? _GEN_8 : temp_result_a; // @[ALU.scala 75:53 ALU.scala 33:30]
  wire [63:0] _GEN_11 = _T_12 & _T_1 ? _GEN_9 : temp_result_b; // @[ALU.scala 75:53 ALU.scala 34:30]
  wire  _GEN_20 = _T_26 & opcode_3 ? io_validin_a : snapshot_valid_a; // @[ALU.scala 103:55 ALU.scala 106:20 ALU.scala 111:20]
  wire  _GEN_24 = opcode_4 & _T_27 ? snapshot_valid_a : _GEN_20; // @[ALU.scala 98:55 ALU.scala 101:20]
  wire  _GEN_28 = ~opcode_4 & ~opcode_3 ? io_validin_a : _GEN_24; // @[ALU.scala 93:49 ALU.scala 96:20]
  wire  _GEN_56 = opcode_8 & opcode_6 & ~opcode_5 ? _GEN_28 : _GEN_28; // @[ALU.scala 114:74]
  wire  gate_valid_a = opcode_8 & ~opcode_6 & opcode_5 ? _GEN_28 : _GEN_56; // @[ALU.scala 92:68]
  wire  _GEN_70 = opcode_0 ? gate_valid_a : temp_valid_a; // @[ALU.scala 181:35 ALU.scala 182:20 ALU.scala 37:29]
  wire  _GEN_72 = ~opcode_0 ? 1'h0 : _GEN_70; // @[ALU.scala 178:29 ALU.scala 179:20]
  assign io_out_a = temp_result_a; // @[ALU.scala 217:12]
  assign io_out_b = temp_result_b; // @[ALU.scala 218:12]
  assign io_validout_a = temp_valid_a; // @[ALU.scala 219:17]
  always @(posedge clock) begin
    if (reset) begin // @[ALU.scala 25:27]
      snapshot_a <= 64'h0; // @[ALU.scala 25:27]
    end else if (opcode_2) begin // @[ALU.scala 160:26]
      snapshot_a <= io_in_a; // @[ALU.scala 161:16]
    end
    if (reset) begin // @[ALU.scala 26:27]
      snapshot_b <= 64'h0; // @[ALU.scala 26:27]
    end else if (opcode_1) begin // @[ALU.scala 168:26]
      snapshot_b <= io_in_b; // @[ALU.scala 169:16]
    end
    if (reset) begin // @[ALU.scala 28:33]
      snapshot_valid_a <= 1'h0; // @[ALU.scala 28:33]
    end else if (opcode_2) begin // @[ALU.scala 160:26]
      snapshot_valid_a <= io_validin_a; // @[ALU.scala 162:22]
    end
    if (reset) begin // @[ALU.scala 33:30]
      temp_result_a <= 64'h0; // @[ALU.scala 33:30]
    end else if (opcode_8 & ~opcode_7) begin // @[ALU.scala 51:47]
      if (opcode_6 & opcode_5) begin // @[ALU.scala 52:49]
        temp_result_a <= _temp_result_a_T_1; // @[ALU.scala 53:21]
      end else begin
        temp_result_a <= _temp_result_a_T; // @[ALU.scala 56:21]
      end
    end else if (opcode_8 & opcode_7) begin // @[ALU.scala 59:53]
      if (_T_5) begin // @[ALU.scala 60:49]
        temp_result_a <= _temp_result_a_T_4; // @[ALU.scala 61:21]
      end else begin
        temp_result_a <= _temp_result_a_T_3; // @[ALU.scala 64:21]
      end
    end else if (~opcode_8 & opcode_7) begin // @[ALU.scala 67:53]
      temp_result_a <= _GEN_4;
    end else begin
      temp_result_a <= _GEN_10;
    end
    if (reset) begin // @[ALU.scala 34:30]
      temp_result_b <= 64'h0; // @[ALU.scala 34:30]
    end else if (opcode_8 & ~opcode_7) begin // @[ALU.scala 51:47]
      temp_result_b <= gate_b;
    end else if (opcode_8 & opcode_7) begin // @[ALU.scala 59:53]
      temp_result_b <= gate_b;
    end else if (~opcode_8 & opcode_7) begin // @[ALU.scala 67:53]
      temp_result_b <= gate_b;
    end else begin
      temp_result_b <= _GEN_11;
    end
    if (reset) begin // @[ALU.scala 37:29]
      temp_valid_a <= 1'h0; // @[ALU.scala 37:29]
    end else if (_T_18) begin // @[ALU.scala 177:47]
      temp_valid_a <= _GEN_72;
    end else begin
      temp_valid_a <= _GEN_72;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  snapshot_a = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  snapshot_b = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  snapshot_valid_a = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  temp_result_a = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  temp_result_b = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  temp_valid_a = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PEcol(
  input          clock,
  input          reset,
  input  [63:0]  io_d_in_0_a,
  input          io_d_in_0_valid_a,
  input  [63:0]  io_d_in_0_b,
  input  [63:0]  io_d_in_1_a,
  input          io_d_in_1_valid_a,
  input  [63:0]  io_d_in_1_b,
  input  [63:0]  io_d_in_2_a,
  input          io_d_in_2_valid_a,
  input  [63:0]  io_d_in_2_b,
  input  [63:0]  io_d_in_3_a,
  input          io_d_in_3_valid_a,
  input  [63:0]  io_d_in_3_b,
  input  [63:0]  io_d_in_4_a,
  input          io_d_in_4_valid_a,
  input  [63:0]  io_d_in_4_b,
  input  [63:0]  io_d_in_5_a,
  input          io_d_in_5_valid_a,
  input  [63:0]  io_d_in_5_b,
  input  [63:0]  io_d_in_6_a,
  input          io_d_in_6_valid_a,
  input  [63:0]  io_d_in_6_b,
  input  [63:0]  io_d_in_7_a,
  input          io_d_in_7_valid_a,
  input  [63:0]  io_d_in_7_b,
  input  [63:0]  io_d_in_8_a,
  input          io_d_in_8_valid_a,
  input  [63:0]  io_d_in_8_b,
  input  [63:0]  io_d_in_9_a,
  input          io_d_in_9_valid_a,
  input  [63:0]  io_d_in_9_b,
  input  [63:0]  io_d_in_10_a,
  input          io_d_in_10_valid_a,
  input  [63:0]  io_d_in_10_b,
  input  [63:0]  io_d_in_11_a,
  input          io_d_in_11_valid_a,
  input  [63:0]  io_d_in_11_b,
  input  [63:0]  io_d_in_12_a,
  input          io_d_in_12_valid_a,
  input  [63:0]  io_d_in_12_b,
  input  [63:0]  io_d_in_13_a,
  input          io_d_in_13_valid_a,
  input  [63:0]  io_d_in_13_b,
  input  [63:0]  io_d_in_14_a,
  input          io_d_in_14_valid_a,
  input  [63:0]  io_d_in_14_b,
  input  [63:0]  io_d_in_15_a,
  input          io_d_in_15_valid_a,
  input  [63:0]  io_d_in_15_b,
  input  [63:0]  io_d_in_16_a,
  input          io_d_in_16_valid_a,
  input  [63:0]  io_d_in_16_b,
  input  [63:0]  io_d_in_17_a,
  input          io_d_in_17_valid_a,
  input  [63:0]  io_d_in_17_b,
  input  [63:0]  io_d_in_18_a,
  input          io_d_in_18_valid_a,
  input  [63:0]  io_d_in_18_b,
  input  [63:0]  io_d_in_19_a,
  input          io_d_in_19_valid_a,
  input  [63:0]  io_d_in_19_b,
  input  [63:0]  io_d_in_20_a,
  input          io_d_in_20_valid_a,
  input  [63:0]  io_d_in_20_b,
  input  [63:0]  io_d_in_21_a,
  input          io_d_in_21_valid_a,
  input  [63:0]  io_d_in_21_b,
  input  [63:0]  io_d_in_22_a,
  input          io_d_in_22_valid_a,
  input  [63:0]  io_d_in_22_b,
  input  [63:0]  io_d_in_23_a,
  input          io_d_in_23_valid_a,
  input  [63:0]  io_d_in_23_b,
  input  [63:0]  io_d_in_24_a,
  input          io_d_in_24_valid_a,
  input  [63:0]  io_d_in_24_b,
  input  [63:0]  io_d_in_25_a,
  input          io_d_in_25_valid_a,
  input  [63:0]  io_d_in_25_b,
  input  [63:0]  io_d_in_26_a,
  input          io_d_in_26_valid_a,
  input  [63:0]  io_d_in_26_b,
  input  [63:0]  io_d_in_27_a,
  input          io_d_in_27_valid_a,
  input  [63:0]  io_d_in_27_b,
  input  [63:0]  io_d_in_28_a,
  input          io_d_in_28_valid_a,
  input  [63:0]  io_d_in_28_b,
  input  [63:0]  io_d_in_29_a,
  input          io_d_in_29_valid_a,
  input  [63:0]  io_d_in_29_b,
  input  [63:0]  io_d_in_30_a,
  input          io_d_in_30_valid_a,
  input  [63:0]  io_d_in_30_b,
  input  [63:0]  io_d_in_31_a,
  input          io_d_in_31_valid_a,
  input  [63:0]  io_d_in_31_b,
  output [63:0]  io_d_out_0_a,
  output         io_d_out_0_valid_a,
  output [63:0]  io_d_out_0_b,
  output [63:0]  io_d_out_1_a,
  output         io_d_out_1_valid_a,
  output [63:0]  io_d_out_1_b,
  output [63:0]  io_d_out_2_a,
  output         io_d_out_2_valid_a,
  output [63:0]  io_d_out_2_b,
  output [63:0]  io_d_out_3_a,
  output         io_d_out_3_valid_a,
  output [63:0]  io_d_out_3_b,
  output [63:0]  io_d_out_4_a,
  output         io_d_out_4_valid_a,
  output [63:0]  io_d_out_4_b,
  output [63:0]  io_d_out_5_a,
  output         io_d_out_5_valid_a,
  output [63:0]  io_d_out_5_b,
  output [63:0]  io_d_out_6_a,
  output         io_d_out_6_valid_a,
  output [63:0]  io_d_out_6_b,
  output [63:0]  io_d_out_7_a,
  output         io_d_out_7_valid_a,
  output [63:0]  io_d_out_7_b,
  output [63:0]  io_d_out_8_a,
  output         io_d_out_8_valid_a,
  output [63:0]  io_d_out_8_b,
  output [63:0]  io_d_out_9_a,
  output         io_d_out_9_valid_a,
  output [63:0]  io_d_out_9_b,
  output [63:0]  io_d_out_10_a,
  output         io_d_out_10_valid_a,
  output [63:0]  io_d_out_10_b,
  output [63:0]  io_d_out_11_a,
  output         io_d_out_11_valid_a,
  output [63:0]  io_d_out_11_b,
  output [63:0]  io_d_out_12_a,
  output         io_d_out_12_valid_a,
  output [63:0]  io_d_out_12_b,
  output [63:0]  io_d_out_13_a,
  output         io_d_out_13_valid_a,
  output [63:0]  io_d_out_13_b,
  output [63:0]  io_d_out_14_a,
  output         io_d_out_14_valid_a,
  output [63:0]  io_d_out_14_b,
  output [63:0]  io_d_out_15_a,
  output         io_d_out_15_valid_a,
  output [63:0]  io_d_out_15_b,
  output [63:0]  io_d_out_16_a,
  output         io_d_out_16_valid_a,
  output [63:0]  io_d_out_16_b,
  output [63:0]  io_d_out_17_a,
  output         io_d_out_17_valid_a,
  output [63:0]  io_d_out_17_b,
  output [63:0]  io_d_out_18_a,
  output         io_d_out_18_valid_a,
  output [63:0]  io_d_out_18_b,
  output [63:0]  io_d_out_19_a,
  output         io_d_out_19_valid_a,
  output [63:0]  io_d_out_19_b,
  output [63:0]  io_d_out_20_a,
  output         io_d_out_20_valid_a,
  output [63:0]  io_d_out_20_b,
  output [63:0]  io_d_out_21_a,
  output         io_d_out_21_valid_a,
  output [63:0]  io_d_out_21_b,
  output [63:0]  io_d_out_22_a,
  output         io_d_out_22_valid_a,
  output [63:0]  io_d_out_22_b,
  output [63:0]  io_d_out_23_a,
  output         io_d_out_23_valid_a,
  output [63:0]  io_d_out_23_b,
  output [63:0]  io_d_out_24_a,
  output         io_d_out_24_valid_a,
  output [63:0]  io_d_out_24_b,
  output [63:0]  io_d_out_25_a,
  output         io_d_out_25_valid_a,
  output [63:0]  io_d_out_25_b,
  output [63:0]  io_d_out_26_a,
  output         io_d_out_26_valid_a,
  output [63:0]  io_d_out_26_b,
  output [63:0]  io_d_out_27_a,
  output         io_d_out_27_valid_a,
  output [63:0]  io_d_out_27_b,
  output [63:0]  io_d_out_28_a,
  output         io_d_out_28_valid_a,
  output [63:0]  io_d_out_28_b,
  output [63:0]  io_d_out_29_a,
  output         io_d_out_29_valid_a,
  output [63:0]  io_d_out_29_b,
  output [63:0]  io_d_out_30_a,
  output         io_d_out_30_valid_a,
  output [63:0]  io_d_out_30_b,
  output [63:0]  io_d_out_31_a,
  output         io_d_out_31_valid_a,
  output [63:0]  io_d_out_31_b,
  input  [1:0]   io_tagin_Tag,
  input  [2:0]   io_tagin_RoundCnt,
  input  [7:0]   io_addrin,
  output [1:0]   io_tagout_Tag,
  output [2:0]   io_tagout_RoundCnt,
  output [7:0]   io_addrout,
  input  [287:0] io_instr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ALU64_32_0_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_0_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_0_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_0_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_0_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_0_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_0_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_0_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_0_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_1_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_1_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_1_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_1_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_1_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_1_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_1_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_1_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_1_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_2_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_2_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_2_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_2_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_2_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_2_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_2_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_2_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_2_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_3_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_3_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_3_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_3_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_3_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_3_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_3_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_3_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_3_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_4_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_4_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_4_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_4_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_4_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_4_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_4_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_4_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_4_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_5_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_5_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_5_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_5_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_5_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_5_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_5_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_5_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_5_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_6_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_6_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_6_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_6_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_6_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_6_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_6_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_6_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_6_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_7_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_7_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_7_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_7_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_7_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_7_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_7_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_7_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_7_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_8_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_8_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_8_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_8_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_8_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_8_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_8_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_8_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_8_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_9_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_9_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_9_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_9_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_9_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_9_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_9_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_9_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_9_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_10_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_10_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_10_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_10_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_10_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_10_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_10_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_10_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_10_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_11_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_11_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_11_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_11_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_11_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_11_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_11_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_11_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_11_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_12_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_12_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_12_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_12_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_12_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_12_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_12_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_12_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_12_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_13_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_13_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_13_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_13_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_13_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_13_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_13_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_13_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_13_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_14_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_14_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_14_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_14_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_14_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_14_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_14_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_14_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_14_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_15_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_15_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_15_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_15_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_15_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_15_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_15_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_15_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_15_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_16_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_16_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_16_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_16_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_16_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_16_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_16_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_16_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_16_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_17_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_17_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_17_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_17_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_17_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_17_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_17_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_17_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_17_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_18_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_18_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_18_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_18_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_18_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_18_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_18_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_18_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_18_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_19_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_19_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_19_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_19_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_19_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_19_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_19_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_19_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_19_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_20_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_20_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_20_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_20_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_20_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_20_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_20_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_20_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_20_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_21_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_21_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_21_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_21_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_21_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_21_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_21_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_21_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_21_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_22_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_22_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_22_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_22_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_22_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_22_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_22_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_22_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_22_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_23_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_23_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_23_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_23_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_23_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_23_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_23_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_23_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_23_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_24_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_24_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_24_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_24_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_24_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_24_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_24_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_24_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_24_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_25_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_25_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_25_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_25_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_25_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_25_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_25_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_25_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_25_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_26_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_26_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_26_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_26_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_26_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_26_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_26_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_26_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_26_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_27_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_27_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_27_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_27_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_27_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_27_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_27_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_27_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_27_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_28_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_28_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_28_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_28_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_28_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_28_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_28_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_28_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_28_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_29_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_29_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_29_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_29_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_29_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_29_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_29_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_29_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_29_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_30_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_30_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_30_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_30_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_30_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_30_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_30_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_30_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_30_io_validout_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_31_clock; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_31_reset; // @[BuildingBlock.scala 231:52]
  wire [8:0] ALU64_32_31_io_opcode; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_31_io_in_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_31_io_in_b; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_31_io_out_a; // @[BuildingBlock.scala 231:52]
  wire [63:0] ALU64_32_31_io_out_b; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_31_io_validin_a; // @[BuildingBlock.scala 231:52]
  wire  ALU64_32_31_io_validout_a; // @[BuildingBlock.scala 231:52]
  reg [1:0] tag_Tag; // @[BuildingBlock.scala 233:20]
  reg [2:0] tag_RoundCnt; // @[BuildingBlock.scala 233:20]
  reg [7:0] addr; // @[BuildingBlock.scala 235:21]
  ALU ALU64_32_0 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_0_clock),
    .reset(ALU64_32_0_reset),
    .io_opcode(ALU64_32_0_io_opcode),
    .io_in_a(ALU64_32_0_io_in_a),
    .io_in_b(ALU64_32_0_io_in_b),
    .io_out_a(ALU64_32_0_io_out_a),
    .io_out_b(ALU64_32_0_io_out_b),
    .io_validin_a(ALU64_32_0_io_validin_a),
    .io_validout_a(ALU64_32_0_io_validout_a)
  );
  ALU ALU64_32_1 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_1_clock),
    .reset(ALU64_32_1_reset),
    .io_opcode(ALU64_32_1_io_opcode),
    .io_in_a(ALU64_32_1_io_in_a),
    .io_in_b(ALU64_32_1_io_in_b),
    .io_out_a(ALU64_32_1_io_out_a),
    .io_out_b(ALU64_32_1_io_out_b),
    .io_validin_a(ALU64_32_1_io_validin_a),
    .io_validout_a(ALU64_32_1_io_validout_a)
  );
  ALU ALU64_32_2 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_2_clock),
    .reset(ALU64_32_2_reset),
    .io_opcode(ALU64_32_2_io_opcode),
    .io_in_a(ALU64_32_2_io_in_a),
    .io_in_b(ALU64_32_2_io_in_b),
    .io_out_a(ALU64_32_2_io_out_a),
    .io_out_b(ALU64_32_2_io_out_b),
    .io_validin_a(ALU64_32_2_io_validin_a),
    .io_validout_a(ALU64_32_2_io_validout_a)
  );
  ALU ALU64_32_3 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_3_clock),
    .reset(ALU64_32_3_reset),
    .io_opcode(ALU64_32_3_io_opcode),
    .io_in_a(ALU64_32_3_io_in_a),
    .io_in_b(ALU64_32_3_io_in_b),
    .io_out_a(ALU64_32_3_io_out_a),
    .io_out_b(ALU64_32_3_io_out_b),
    .io_validin_a(ALU64_32_3_io_validin_a),
    .io_validout_a(ALU64_32_3_io_validout_a)
  );
  ALU ALU64_32_4 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_4_clock),
    .reset(ALU64_32_4_reset),
    .io_opcode(ALU64_32_4_io_opcode),
    .io_in_a(ALU64_32_4_io_in_a),
    .io_in_b(ALU64_32_4_io_in_b),
    .io_out_a(ALU64_32_4_io_out_a),
    .io_out_b(ALU64_32_4_io_out_b),
    .io_validin_a(ALU64_32_4_io_validin_a),
    .io_validout_a(ALU64_32_4_io_validout_a)
  );
  ALU ALU64_32_5 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_5_clock),
    .reset(ALU64_32_5_reset),
    .io_opcode(ALU64_32_5_io_opcode),
    .io_in_a(ALU64_32_5_io_in_a),
    .io_in_b(ALU64_32_5_io_in_b),
    .io_out_a(ALU64_32_5_io_out_a),
    .io_out_b(ALU64_32_5_io_out_b),
    .io_validin_a(ALU64_32_5_io_validin_a),
    .io_validout_a(ALU64_32_5_io_validout_a)
  );
  ALU ALU64_32_6 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_6_clock),
    .reset(ALU64_32_6_reset),
    .io_opcode(ALU64_32_6_io_opcode),
    .io_in_a(ALU64_32_6_io_in_a),
    .io_in_b(ALU64_32_6_io_in_b),
    .io_out_a(ALU64_32_6_io_out_a),
    .io_out_b(ALU64_32_6_io_out_b),
    .io_validin_a(ALU64_32_6_io_validin_a),
    .io_validout_a(ALU64_32_6_io_validout_a)
  );
  ALU ALU64_32_7 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_7_clock),
    .reset(ALU64_32_7_reset),
    .io_opcode(ALU64_32_7_io_opcode),
    .io_in_a(ALU64_32_7_io_in_a),
    .io_in_b(ALU64_32_7_io_in_b),
    .io_out_a(ALU64_32_7_io_out_a),
    .io_out_b(ALU64_32_7_io_out_b),
    .io_validin_a(ALU64_32_7_io_validin_a),
    .io_validout_a(ALU64_32_7_io_validout_a)
  );
  ALU ALU64_32_8 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_8_clock),
    .reset(ALU64_32_8_reset),
    .io_opcode(ALU64_32_8_io_opcode),
    .io_in_a(ALU64_32_8_io_in_a),
    .io_in_b(ALU64_32_8_io_in_b),
    .io_out_a(ALU64_32_8_io_out_a),
    .io_out_b(ALU64_32_8_io_out_b),
    .io_validin_a(ALU64_32_8_io_validin_a),
    .io_validout_a(ALU64_32_8_io_validout_a)
  );
  ALU ALU64_32_9 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_9_clock),
    .reset(ALU64_32_9_reset),
    .io_opcode(ALU64_32_9_io_opcode),
    .io_in_a(ALU64_32_9_io_in_a),
    .io_in_b(ALU64_32_9_io_in_b),
    .io_out_a(ALU64_32_9_io_out_a),
    .io_out_b(ALU64_32_9_io_out_b),
    .io_validin_a(ALU64_32_9_io_validin_a),
    .io_validout_a(ALU64_32_9_io_validout_a)
  );
  ALU ALU64_32_10 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_10_clock),
    .reset(ALU64_32_10_reset),
    .io_opcode(ALU64_32_10_io_opcode),
    .io_in_a(ALU64_32_10_io_in_a),
    .io_in_b(ALU64_32_10_io_in_b),
    .io_out_a(ALU64_32_10_io_out_a),
    .io_out_b(ALU64_32_10_io_out_b),
    .io_validin_a(ALU64_32_10_io_validin_a),
    .io_validout_a(ALU64_32_10_io_validout_a)
  );
  ALU ALU64_32_11 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_11_clock),
    .reset(ALU64_32_11_reset),
    .io_opcode(ALU64_32_11_io_opcode),
    .io_in_a(ALU64_32_11_io_in_a),
    .io_in_b(ALU64_32_11_io_in_b),
    .io_out_a(ALU64_32_11_io_out_a),
    .io_out_b(ALU64_32_11_io_out_b),
    .io_validin_a(ALU64_32_11_io_validin_a),
    .io_validout_a(ALU64_32_11_io_validout_a)
  );
  ALU ALU64_32_12 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_12_clock),
    .reset(ALU64_32_12_reset),
    .io_opcode(ALU64_32_12_io_opcode),
    .io_in_a(ALU64_32_12_io_in_a),
    .io_in_b(ALU64_32_12_io_in_b),
    .io_out_a(ALU64_32_12_io_out_a),
    .io_out_b(ALU64_32_12_io_out_b),
    .io_validin_a(ALU64_32_12_io_validin_a),
    .io_validout_a(ALU64_32_12_io_validout_a)
  );
  ALU ALU64_32_13 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_13_clock),
    .reset(ALU64_32_13_reset),
    .io_opcode(ALU64_32_13_io_opcode),
    .io_in_a(ALU64_32_13_io_in_a),
    .io_in_b(ALU64_32_13_io_in_b),
    .io_out_a(ALU64_32_13_io_out_a),
    .io_out_b(ALU64_32_13_io_out_b),
    .io_validin_a(ALU64_32_13_io_validin_a),
    .io_validout_a(ALU64_32_13_io_validout_a)
  );
  ALU ALU64_32_14 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_14_clock),
    .reset(ALU64_32_14_reset),
    .io_opcode(ALU64_32_14_io_opcode),
    .io_in_a(ALU64_32_14_io_in_a),
    .io_in_b(ALU64_32_14_io_in_b),
    .io_out_a(ALU64_32_14_io_out_a),
    .io_out_b(ALU64_32_14_io_out_b),
    .io_validin_a(ALU64_32_14_io_validin_a),
    .io_validout_a(ALU64_32_14_io_validout_a)
  );
  ALU ALU64_32_15 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_15_clock),
    .reset(ALU64_32_15_reset),
    .io_opcode(ALU64_32_15_io_opcode),
    .io_in_a(ALU64_32_15_io_in_a),
    .io_in_b(ALU64_32_15_io_in_b),
    .io_out_a(ALU64_32_15_io_out_a),
    .io_out_b(ALU64_32_15_io_out_b),
    .io_validin_a(ALU64_32_15_io_validin_a),
    .io_validout_a(ALU64_32_15_io_validout_a)
  );
  ALU ALU64_32_16 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_16_clock),
    .reset(ALU64_32_16_reset),
    .io_opcode(ALU64_32_16_io_opcode),
    .io_in_a(ALU64_32_16_io_in_a),
    .io_in_b(ALU64_32_16_io_in_b),
    .io_out_a(ALU64_32_16_io_out_a),
    .io_out_b(ALU64_32_16_io_out_b),
    .io_validin_a(ALU64_32_16_io_validin_a),
    .io_validout_a(ALU64_32_16_io_validout_a)
  );
  ALU ALU64_32_17 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_17_clock),
    .reset(ALU64_32_17_reset),
    .io_opcode(ALU64_32_17_io_opcode),
    .io_in_a(ALU64_32_17_io_in_a),
    .io_in_b(ALU64_32_17_io_in_b),
    .io_out_a(ALU64_32_17_io_out_a),
    .io_out_b(ALU64_32_17_io_out_b),
    .io_validin_a(ALU64_32_17_io_validin_a),
    .io_validout_a(ALU64_32_17_io_validout_a)
  );
  ALU ALU64_32_18 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_18_clock),
    .reset(ALU64_32_18_reset),
    .io_opcode(ALU64_32_18_io_opcode),
    .io_in_a(ALU64_32_18_io_in_a),
    .io_in_b(ALU64_32_18_io_in_b),
    .io_out_a(ALU64_32_18_io_out_a),
    .io_out_b(ALU64_32_18_io_out_b),
    .io_validin_a(ALU64_32_18_io_validin_a),
    .io_validout_a(ALU64_32_18_io_validout_a)
  );
  ALU ALU64_32_19 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_19_clock),
    .reset(ALU64_32_19_reset),
    .io_opcode(ALU64_32_19_io_opcode),
    .io_in_a(ALU64_32_19_io_in_a),
    .io_in_b(ALU64_32_19_io_in_b),
    .io_out_a(ALU64_32_19_io_out_a),
    .io_out_b(ALU64_32_19_io_out_b),
    .io_validin_a(ALU64_32_19_io_validin_a),
    .io_validout_a(ALU64_32_19_io_validout_a)
  );
  ALU ALU64_32_20 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_20_clock),
    .reset(ALU64_32_20_reset),
    .io_opcode(ALU64_32_20_io_opcode),
    .io_in_a(ALU64_32_20_io_in_a),
    .io_in_b(ALU64_32_20_io_in_b),
    .io_out_a(ALU64_32_20_io_out_a),
    .io_out_b(ALU64_32_20_io_out_b),
    .io_validin_a(ALU64_32_20_io_validin_a),
    .io_validout_a(ALU64_32_20_io_validout_a)
  );
  ALU ALU64_32_21 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_21_clock),
    .reset(ALU64_32_21_reset),
    .io_opcode(ALU64_32_21_io_opcode),
    .io_in_a(ALU64_32_21_io_in_a),
    .io_in_b(ALU64_32_21_io_in_b),
    .io_out_a(ALU64_32_21_io_out_a),
    .io_out_b(ALU64_32_21_io_out_b),
    .io_validin_a(ALU64_32_21_io_validin_a),
    .io_validout_a(ALU64_32_21_io_validout_a)
  );
  ALU ALU64_32_22 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_22_clock),
    .reset(ALU64_32_22_reset),
    .io_opcode(ALU64_32_22_io_opcode),
    .io_in_a(ALU64_32_22_io_in_a),
    .io_in_b(ALU64_32_22_io_in_b),
    .io_out_a(ALU64_32_22_io_out_a),
    .io_out_b(ALU64_32_22_io_out_b),
    .io_validin_a(ALU64_32_22_io_validin_a),
    .io_validout_a(ALU64_32_22_io_validout_a)
  );
  ALU ALU64_32_23 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_23_clock),
    .reset(ALU64_32_23_reset),
    .io_opcode(ALU64_32_23_io_opcode),
    .io_in_a(ALU64_32_23_io_in_a),
    .io_in_b(ALU64_32_23_io_in_b),
    .io_out_a(ALU64_32_23_io_out_a),
    .io_out_b(ALU64_32_23_io_out_b),
    .io_validin_a(ALU64_32_23_io_validin_a),
    .io_validout_a(ALU64_32_23_io_validout_a)
  );
  ALU ALU64_32_24 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_24_clock),
    .reset(ALU64_32_24_reset),
    .io_opcode(ALU64_32_24_io_opcode),
    .io_in_a(ALU64_32_24_io_in_a),
    .io_in_b(ALU64_32_24_io_in_b),
    .io_out_a(ALU64_32_24_io_out_a),
    .io_out_b(ALU64_32_24_io_out_b),
    .io_validin_a(ALU64_32_24_io_validin_a),
    .io_validout_a(ALU64_32_24_io_validout_a)
  );
  ALU ALU64_32_25 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_25_clock),
    .reset(ALU64_32_25_reset),
    .io_opcode(ALU64_32_25_io_opcode),
    .io_in_a(ALU64_32_25_io_in_a),
    .io_in_b(ALU64_32_25_io_in_b),
    .io_out_a(ALU64_32_25_io_out_a),
    .io_out_b(ALU64_32_25_io_out_b),
    .io_validin_a(ALU64_32_25_io_validin_a),
    .io_validout_a(ALU64_32_25_io_validout_a)
  );
  ALU ALU64_32_26 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_26_clock),
    .reset(ALU64_32_26_reset),
    .io_opcode(ALU64_32_26_io_opcode),
    .io_in_a(ALU64_32_26_io_in_a),
    .io_in_b(ALU64_32_26_io_in_b),
    .io_out_a(ALU64_32_26_io_out_a),
    .io_out_b(ALU64_32_26_io_out_b),
    .io_validin_a(ALU64_32_26_io_validin_a),
    .io_validout_a(ALU64_32_26_io_validout_a)
  );
  ALU ALU64_32_27 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_27_clock),
    .reset(ALU64_32_27_reset),
    .io_opcode(ALU64_32_27_io_opcode),
    .io_in_a(ALU64_32_27_io_in_a),
    .io_in_b(ALU64_32_27_io_in_b),
    .io_out_a(ALU64_32_27_io_out_a),
    .io_out_b(ALU64_32_27_io_out_b),
    .io_validin_a(ALU64_32_27_io_validin_a),
    .io_validout_a(ALU64_32_27_io_validout_a)
  );
  ALU ALU64_32_28 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_28_clock),
    .reset(ALU64_32_28_reset),
    .io_opcode(ALU64_32_28_io_opcode),
    .io_in_a(ALU64_32_28_io_in_a),
    .io_in_b(ALU64_32_28_io_in_b),
    .io_out_a(ALU64_32_28_io_out_a),
    .io_out_b(ALU64_32_28_io_out_b),
    .io_validin_a(ALU64_32_28_io_validin_a),
    .io_validout_a(ALU64_32_28_io_validout_a)
  );
  ALU ALU64_32_29 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_29_clock),
    .reset(ALU64_32_29_reset),
    .io_opcode(ALU64_32_29_io_opcode),
    .io_in_a(ALU64_32_29_io_in_a),
    .io_in_b(ALU64_32_29_io_in_b),
    .io_out_a(ALU64_32_29_io_out_a),
    .io_out_b(ALU64_32_29_io_out_b),
    .io_validin_a(ALU64_32_29_io_validin_a),
    .io_validout_a(ALU64_32_29_io_validout_a)
  );
  ALU ALU64_32_30 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_30_clock),
    .reset(ALU64_32_30_reset),
    .io_opcode(ALU64_32_30_io_opcode),
    .io_in_a(ALU64_32_30_io_in_a),
    .io_in_b(ALU64_32_30_io_in_b),
    .io_out_a(ALU64_32_30_io_out_a),
    .io_out_b(ALU64_32_30_io_out_b),
    .io_validin_a(ALU64_32_30_io_validin_a),
    .io_validout_a(ALU64_32_30_io_validout_a)
  );
  ALU ALU64_32_31 ( // @[BuildingBlock.scala 231:52]
    .clock(ALU64_32_31_clock),
    .reset(ALU64_32_31_reset),
    .io_opcode(ALU64_32_31_io_opcode),
    .io_in_a(ALU64_32_31_io_in_a),
    .io_in_b(ALU64_32_31_io_in_b),
    .io_out_a(ALU64_32_31_io_out_a),
    .io_out_b(ALU64_32_31_io_out_b),
    .io_validin_a(ALU64_32_31_io_validin_a),
    .io_validout_a(ALU64_32_31_io_validout_a)
  );
  assign io_d_out_0_a = ALU64_32_0_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_0_valid_a = ALU64_32_0_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_0_b = ALU64_32_0_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_1_a = ALU64_32_1_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_1_valid_a = ALU64_32_1_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_1_b = ALU64_32_1_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_2_a = ALU64_32_2_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_2_valid_a = ALU64_32_2_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_2_b = ALU64_32_2_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_3_a = ALU64_32_3_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_3_valid_a = ALU64_32_3_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_3_b = ALU64_32_3_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_4_a = ALU64_32_4_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_4_valid_a = ALU64_32_4_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_4_b = ALU64_32_4_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_5_a = ALU64_32_5_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_5_valid_a = ALU64_32_5_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_5_b = ALU64_32_5_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_6_a = ALU64_32_6_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_6_valid_a = ALU64_32_6_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_6_b = ALU64_32_6_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_7_a = ALU64_32_7_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_7_valid_a = ALU64_32_7_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_7_b = ALU64_32_7_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_8_a = ALU64_32_8_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_8_valid_a = ALU64_32_8_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_8_b = ALU64_32_8_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_9_a = ALU64_32_9_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_9_valid_a = ALU64_32_9_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_9_b = ALU64_32_9_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_10_a = ALU64_32_10_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_10_valid_a = ALU64_32_10_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_10_b = ALU64_32_10_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_11_a = ALU64_32_11_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_11_valid_a = ALU64_32_11_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_11_b = ALU64_32_11_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_12_a = ALU64_32_12_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_12_valid_a = ALU64_32_12_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_12_b = ALU64_32_12_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_13_a = ALU64_32_13_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_13_valid_a = ALU64_32_13_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_13_b = ALU64_32_13_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_14_a = ALU64_32_14_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_14_valid_a = ALU64_32_14_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_14_b = ALU64_32_14_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_15_a = ALU64_32_15_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_15_valid_a = ALU64_32_15_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_15_b = ALU64_32_15_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_16_a = ALU64_32_16_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_16_valid_a = ALU64_32_16_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_16_b = ALU64_32_16_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_17_a = ALU64_32_17_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_17_valid_a = ALU64_32_17_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_17_b = ALU64_32_17_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_18_a = ALU64_32_18_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_18_valid_a = ALU64_32_18_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_18_b = ALU64_32_18_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_19_a = ALU64_32_19_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_19_valid_a = ALU64_32_19_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_19_b = ALU64_32_19_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_20_a = ALU64_32_20_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_20_valid_a = ALU64_32_20_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_20_b = ALU64_32_20_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_21_a = ALU64_32_21_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_21_valid_a = ALU64_32_21_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_21_b = ALU64_32_21_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_22_a = ALU64_32_22_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_22_valid_a = ALU64_32_22_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_22_b = ALU64_32_22_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_23_a = ALU64_32_23_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_23_valid_a = ALU64_32_23_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_23_b = ALU64_32_23_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_24_a = ALU64_32_24_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_24_valid_a = ALU64_32_24_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_24_b = ALU64_32_24_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_25_a = ALU64_32_25_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_25_valid_a = ALU64_32_25_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_25_b = ALU64_32_25_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_26_a = ALU64_32_26_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_26_valid_a = ALU64_32_26_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_26_b = ALU64_32_26_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_27_a = ALU64_32_27_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_27_valid_a = ALU64_32_27_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_27_b = ALU64_32_27_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_28_a = ALU64_32_28_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_28_valid_a = ALU64_32_28_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_28_b = ALU64_32_28_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_29_a = ALU64_32_29_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_29_valid_a = ALU64_32_29_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_29_b = ALU64_32_29_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_30_a = ALU64_32_30_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_30_valid_a = ALU64_32_30_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_30_b = ALU64_32_30_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_d_out_31_a = ALU64_32_31_io_out_a; // @[BuildingBlock.scala 249:19]
  assign io_d_out_31_valid_a = ALU64_32_31_io_validout_a; // @[BuildingBlock.scala 251:25]
  assign io_d_out_31_b = ALU64_32_31_io_out_b; // @[BuildingBlock.scala 250:19]
  assign io_tagout_Tag = tag_Tag; // @[BuildingBlock.scala 234:13]
  assign io_tagout_RoundCnt = tag_RoundCnt; // @[BuildingBlock.scala 234:13]
  assign io_addrout = addr; // @[BuildingBlock.scala 236:14]
  assign ALU64_32_0_clock = clock;
  assign ALU64_32_0_reset = reset;
  assign ALU64_32_0_io_opcode = io_instr[287:279]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_0_io_in_a = io_d_in_0_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_0_io_in_b = io_d_in_0_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_0_io_validin_a = io_d_in_0_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_1_clock = clock;
  assign ALU64_32_1_reset = reset;
  assign ALU64_32_1_io_opcode = io_instr[278:270]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_1_io_in_a = io_d_in_1_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_1_io_in_b = io_d_in_1_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_1_io_validin_a = io_d_in_1_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_2_clock = clock;
  assign ALU64_32_2_reset = reset;
  assign ALU64_32_2_io_opcode = io_instr[269:261]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_2_io_in_a = io_d_in_2_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_2_io_in_b = io_d_in_2_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_2_io_validin_a = io_d_in_2_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_3_clock = clock;
  assign ALU64_32_3_reset = reset;
  assign ALU64_32_3_io_opcode = io_instr[260:252]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_3_io_in_a = io_d_in_3_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_3_io_in_b = io_d_in_3_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_3_io_validin_a = io_d_in_3_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_4_clock = clock;
  assign ALU64_32_4_reset = reset;
  assign ALU64_32_4_io_opcode = io_instr[251:243]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_4_io_in_a = io_d_in_4_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_4_io_in_b = io_d_in_4_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_4_io_validin_a = io_d_in_4_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_5_clock = clock;
  assign ALU64_32_5_reset = reset;
  assign ALU64_32_5_io_opcode = io_instr[242:234]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_5_io_in_a = io_d_in_5_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_5_io_in_b = io_d_in_5_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_5_io_validin_a = io_d_in_5_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_6_clock = clock;
  assign ALU64_32_6_reset = reset;
  assign ALU64_32_6_io_opcode = io_instr[233:225]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_6_io_in_a = io_d_in_6_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_6_io_in_b = io_d_in_6_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_6_io_validin_a = io_d_in_6_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_7_clock = clock;
  assign ALU64_32_7_reset = reset;
  assign ALU64_32_7_io_opcode = io_instr[224:216]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_7_io_in_a = io_d_in_7_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_7_io_in_b = io_d_in_7_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_7_io_validin_a = io_d_in_7_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_8_clock = clock;
  assign ALU64_32_8_reset = reset;
  assign ALU64_32_8_io_opcode = io_instr[215:207]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_8_io_in_a = io_d_in_8_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_8_io_in_b = io_d_in_8_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_8_io_validin_a = io_d_in_8_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_9_clock = clock;
  assign ALU64_32_9_reset = reset;
  assign ALU64_32_9_io_opcode = io_instr[206:198]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_9_io_in_a = io_d_in_9_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_9_io_in_b = io_d_in_9_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_9_io_validin_a = io_d_in_9_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_10_clock = clock;
  assign ALU64_32_10_reset = reset;
  assign ALU64_32_10_io_opcode = io_instr[197:189]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_10_io_in_a = io_d_in_10_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_10_io_in_b = io_d_in_10_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_10_io_validin_a = io_d_in_10_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_11_clock = clock;
  assign ALU64_32_11_reset = reset;
  assign ALU64_32_11_io_opcode = io_instr[188:180]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_11_io_in_a = io_d_in_11_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_11_io_in_b = io_d_in_11_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_11_io_validin_a = io_d_in_11_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_12_clock = clock;
  assign ALU64_32_12_reset = reset;
  assign ALU64_32_12_io_opcode = io_instr[179:171]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_12_io_in_a = io_d_in_12_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_12_io_in_b = io_d_in_12_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_12_io_validin_a = io_d_in_12_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_13_clock = clock;
  assign ALU64_32_13_reset = reset;
  assign ALU64_32_13_io_opcode = io_instr[170:162]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_13_io_in_a = io_d_in_13_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_13_io_in_b = io_d_in_13_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_13_io_validin_a = io_d_in_13_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_14_clock = clock;
  assign ALU64_32_14_reset = reset;
  assign ALU64_32_14_io_opcode = io_instr[161:153]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_14_io_in_a = io_d_in_14_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_14_io_in_b = io_d_in_14_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_14_io_validin_a = io_d_in_14_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_15_clock = clock;
  assign ALU64_32_15_reset = reset;
  assign ALU64_32_15_io_opcode = io_instr[152:144]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_15_io_in_a = io_d_in_15_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_15_io_in_b = io_d_in_15_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_15_io_validin_a = io_d_in_15_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_16_clock = clock;
  assign ALU64_32_16_reset = reset;
  assign ALU64_32_16_io_opcode = io_instr[143:135]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_16_io_in_a = io_d_in_16_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_16_io_in_b = io_d_in_16_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_16_io_validin_a = io_d_in_16_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_17_clock = clock;
  assign ALU64_32_17_reset = reset;
  assign ALU64_32_17_io_opcode = io_instr[134:126]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_17_io_in_a = io_d_in_17_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_17_io_in_b = io_d_in_17_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_17_io_validin_a = io_d_in_17_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_18_clock = clock;
  assign ALU64_32_18_reset = reset;
  assign ALU64_32_18_io_opcode = io_instr[125:117]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_18_io_in_a = io_d_in_18_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_18_io_in_b = io_d_in_18_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_18_io_validin_a = io_d_in_18_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_19_clock = clock;
  assign ALU64_32_19_reset = reset;
  assign ALU64_32_19_io_opcode = io_instr[116:108]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_19_io_in_a = io_d_in_19_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_19_io_in_b = io_d_in_19_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_19_io_validin_a = io_d_in_19_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_20_clock = clock;
  assign ALU64_32_20_reset = reset;
  assign ALU64_32_20_io_opcode = io_instr[107:99]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_20_io_in_a = io_d_in_20_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_20_io_in_b = io_d_in_20_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_20_io_validin_a = io_d_in_20_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_21_clock = clock;
  assign ALU64_32_21_reset = reset;
  assign ALU64_32_21_io_opcode = io_instr[98:90]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_21_io_in_a = io_d_in_21_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_21_io_in_b = io_d_in_21_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_21_io_validin_a = io_d_in_21_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_22_clock = clock;
  assign ALU64_32_22_reset = reset;
  assign ALU64_32_22_io_opcode = io_instr[89:81]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_22_io_in_a = io_d_in_22_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_22_io_in_b = io_d_in_22_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_22_io_validin_a = io_d_in_22_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_23_clock = clock;
  assign ALU64_32_23_reset = reset;
  assign ALU64_32_23_io_opcode = io_instr[80:72]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_23_io_in_a = io_d_in_23_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_23_io_in_b = io_d_in_23_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_23_io_validin_a = io_d_in_23_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_24_clock = clock;
  assign ALU64_32_24_reset = reset;
  assign ALU64_32_24_io_opcode = io_instr[71:63]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_24_io_in_a = io_d_in_24_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_24_io_in_b = io_d_in_24_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_24_io_validin_a = io_d_in_24_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_25_clock = clock;
  assign ALU64_32_25_reset = reset;
  assign ALU64_32_25_io_opcode = io_instr[62:54]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_25_io_in_a = io_d_in_25_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_25_io_in_b = io_d_in_25_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_25_io_validin_a = io_d_in_25_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_26_clock = clock;
  assign ALU64_32_26_reset = reset;
  assign ALU64_32_26_io_opcode = io_instr[53:45]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_26_io_in_a = io_d_in_26_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_26_io_in_b = io_d_in_26_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_26_io_validin_a = io_d_in_26_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_27_clock = clock;
  assign ALU64_32_27_reset = reset;
  assign ALU64_32_27_io_opcode = io_instr[44:36]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_27_io_in_a = io_d_in_27_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_27_io_in_b = io_d_in_27_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_27_io_validin_a = io_d_in_27_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_28_clock = clock;
  assign ALU64_32_28_reset = reset;
  assign ALU64_32_28_io_opcode = io_instr[35:27]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_28_io_in_a = io_d_in_28_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_28_io_in_b = io_d_in_28_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_28_io_validin_a = io_d_in_28_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_29_clock = clock;
  assign ALU64_32_29_reset = reset;
  assign ALU64_32_29_io_opcode = io_instr[26:18]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_29_io_in_a = io_d_in_29_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_29_io_in_b = io_d_in_29_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_29_io_validin_a = io_d_in_29_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_30_clock = clock;
  assign ALU64_32_30_reset = reset;
  assign ALU64_32_30_io_opcode = io_instr[17:9]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_30_io_in_a = io_d_in_30_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_30_io_in_b = io_d_in_30_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_30_io_validin_a = io_d_in_30_valid_a; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_31_clock = clock;
  assign ALU64_32_31_reset = reset;
  assign ALU64_32_31_io_opcode = io_instr[8:0]; // @[BuildingBlock.scala 245:38]
  assign ALU64_32_31_io_in_a = io_d_in_31_a; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_31_io_in_b = io_d_in_31_b; // @[BuildingBlock.scala 242:25]
  assign ALU64_32_31_io_validin_a = io_d_in_31_valid_a; // @[BuildingBlock.scala 243:30]
  always @(posedge clock) begin
    tag_Tag <= io_tagin_Tag; // @[BuildingBlock.scala 233:20]
    tag_RoundCnt <= io_tagin_RoundCnt; // @[BuildingBlock.scala 233:20]
    addr <= io_addrin; // @[BuildingBlock.scala 235:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_Tag = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  tag_RoundCnt = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  addr = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CrossBarCell(
  input  [64:0] io_fw_left,
  input  [64:0] io_fw_top,
  output [64:0] io_fw_bottom,
  output [64:0] io_fw_right,
  input         io_sel
);
  assign io_fw_bottom = io_sel ? io_fw_left : io_fw_top; // @[CrossBarSwitch.scala 16:17 CrossBarSwitch.scala 17:18 CrossBarSwitch.scala 19:18]
  assign io_fw_right = io_fw_left; // @[CrossBarSwitch.scala 15:15]
endmodule
module CrossBarSwitch(
  input         clock,
  input  [64:0] io_fw_left_0,
  input  [64:0] io_fw_left_1,
  input  [64:0] io_fw_left_2,
  input  [64:0] io_fw_left_3,
  output [64:0] io_fw_bottom_0,
  output [64:0] io_fw_bottom_1,
  output [64:0] io_fw_bottom_2,
  output [64:0] io_fw_bottom_3,
  input  [1:0]  io_select_0,
  input  [1:0]  io_select_1,
  input  [1:0]  io_select_2,
  input  [1:0]  io_select_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [95:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [64:0] cells_2d_0_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_0_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_0_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_0_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_0_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_1_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_1_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_1_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_1_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_1_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_2_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_2_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_2_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_2_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_2_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_3_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_3_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_3_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_3_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_3_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_4_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_4_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_4_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_4_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_4_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_5_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_5_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_5_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_5_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_5_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_6_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_6_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_6_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_6_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_6_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_7_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_7_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_7_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_7_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_7_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_8_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_8_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_8_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_8_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_8_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_9_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_9_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_9_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_9_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_9_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_10_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_10_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_10_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_10_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_10_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_11_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_11_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_11_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_11_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_11_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_12_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_12_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_12_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_12_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_12_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_13_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_13_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_13_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_13_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_13_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_14_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_14_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_14_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_14_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_14_io_sel; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_15_io_fw_left; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_15_io_fw_top; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_15_io_fw_bottom; // @[CrossBarSwitch.scala 100:53]
  wire [64:0] cells_2d_15_io_fw_right; // @[CrossBarSwitch.scala 100:53]
  wire  cells_2d_15_io_sel; // @[CrossBarSwitch.scala 100:53]
  reg [64:0] fw_bottom_reg_0; // @[CrossBarSwitch.scala 97:26]
  reg [64:0] fw_bottom_reg_1; // @[CrossBarSwitch.scala 97:26]
  reg [64:0] fw_bottom_reg_2; // @[CrossBarSwitch.scala 97:26]
  reg [64:0] fw_bottom_reg_3; // @[CrossBarSwitch.scala 97:26]
  wire [3:0] select_onehot_0 = 4'h1 << io_select_0; // @[OneHot.scala 65:12]
  wire [3:0] select_onehot_1 = 4'h1 << io_select_1; // @[OneHot.scala 65:12]
  wire [3:0] select_onehot_2 = 4'h1 << io_select_2; // @[OneHot.scala 65:12]
  wire [3:0] select_onehot_3 = 4'h1 << io_select_3; // @[OneHot.scala 65:12]
  CrossBarCell cells_2d_0 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_0_io_fw_left),
    .io_fw_top(cells_2d_0_io_fw_top),
    .io_fw_bottom(cells_2d_0_io_fw_bottom),
    .io_fw_right(cells_2d_0_io_fw_right),
    .io_sel(cells_2d_0_io_sel)
  );
  CrossBarCell cells_2d_1 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_1_io_fw_left),
    .io_fw_top(cells_2d_1_io_fw_top),
    .io_fw_bottom(cells_2d_1_io_fw_bottom),
    .io_fw_right(cells_2d_1_io_fw_right),
    .io_sel(cells_2d_1_io_sel)
  );
  CrossBarCell cells_2d_2 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_2_io_fw_left),
    .io_fw_top(cells_2d_2_io_fw_top),
    .io_fw_bottom(cells_2d_2_io_fw_bottom),
    .io_fw_right(cells_2d_2_io_fw_right),
    .io_sel(cells_2d_2_io_sel)
  );
  CrossBarCell cells_2d_3 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_3_io_fw_left),
    .io_fw_top(cells_2d_3_io_fw_top),
    .io_fw_bottom(cells_2d_3_io_fw_bottom),
    .io_fw_right(cells_2d_3_io_fw_right),
    .io_sel(cells_2d_3_io_sel)
  );
  CrossBarCell cells_2d_4 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_4_io_fw_left),
    .io_fw_top(cells_2d_4_io_fw_top),
    .io_fw_bottom(cells_2d_4_io_fw_bottom),
    .io_fw_right(cells_2d_4_io_fw_right),
    .io_sel(cells_2d_4_io_sel)
  );
  CrossBarCell cells_2d_5 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_5_io_fw_left),
    .io_fw_top(cells_2d_5_io_fw_top),
    .io_fw_bottom(cells_2d_5_io_fw_bottom),
    .io_fw_right(cells_2d_5_io_fw_right),
    .io_sel(cells_2d_5_io_sel)
  );
  CrossBarCell cells_2d_6 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_6_io_fw_left),
    .io_fw_top(cells_2d_6_io_fw_top),
    .io_fw_bottom(cells_2d_6_io_fw_bottom),
    .io_fw_right(cells_2d_6_io_fw_right),
    .io_sel(cells_2d_6_io_sel)
  );
  CrossBarCell cells_2d_7 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_7_io_fw_left),
    .io_fw_top(cells_2d_7_io_fw_top),
    .io_fw_bottom(cells_2d_7_io_fw_bottom),
    .io_fw_right(cells_2d_7_io_fw_right),
    .io_sel(cells_2d_7_io_sel)
  );
  CrossBarCell cells_2d_8 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_8_io_fw_left),
    .io_fw_top(cells_2d_8_io_fw_top),
    .io_fw_bottom(cells_2d_8_io_fw_bottom),
    .io_fw_right(cells_2d_8_io_fw_right),
    .io_sel(cells_2d_8_io_sel)
  );
  CrossBarCell cells_2d_9 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_9_io_fw_left),
    .io_fw_top(cells_2d_9_io_fw_top),
    .io_fw_bottom(cells_2d_9_io_fw_bottom),
    .io_fw_right(cells_2d_9_io_fw_right),
    .io_sel(cells_2d_9_io_sel)
  );
  CrossBarCell cells_2d_10 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_10_io_fw_left),
    .io_fw_top(cells_2d_10_io_fw_top),
    .io_fw_bottom(cells_2d_10_io_fw_bottom),
    .io_fw_right(cells_2d_10_io_fw_right),
    .io_sel(cells_2d_10_io_sel)
  );
  CrossBarCell cells_2d_11 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_11_io_fw_left),
    .io_fw_top(cells_2d_11_io_fw_top),
    .io_fw_bottom(cells_2d_11_io_fw_bottom),
    .io_fw_right(cells_2d_11_io_fw_right),
    .io_sel(cells_2d_11_io_sel)
  );
  CrossBarCell cells_2d_12 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_12_io_fw_left),
    .io_fw_top(cells_2d_12_io_fw_top),
    .io_fw_bottom(cells_2d_12_io_fw_bottom),
    .io_fw_right(cells_2d_12_io_fw_right),
    .io_sel(cells_2d_12_io_sel)
  );
  CrossBarCell cells_2d_13 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_13_io_fw_left),
    .io_fw_top(cells_2d_13_io_fw_top),
    .io_fw_bottom(cells_2d_13_io_fw_bottom),
    .io_fw_right(cells_2d_13_io_fw_right),
    .io_sel(cells_2d_13_io_sel)
  );
  CrossBarCell cells_2d_14 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_14_io_fw_left),
    .io_fw_top(cells_2d_14_io_fw_top),
    .io_fw_bottom(cells_2d_14_io_fw_bottom),
    .io_fw_right(cells_2d_14_io_fw_right),
    .io_sel(cells_2d_14_io_sel)
  );
  CrossBarCell cells_2d_15 ( // @[CrossBarSwitch.scala 100:53]
    .io_fw_left(cells_2d_15_io_fw_left),
    .io_fw_top(cells_2d_15_io_fw_top),
    .io_fw_bottom(cells_2d_15_io_fw_bottom),
    .io_fw_right(cells_2d_15_io_fw_right),
    .io_sel(cells_2d_15_io_sel)
  );
  assign io_fw_bottom_0 = fw_bottom_reg_0; // @[CrossBarSwitch.scala 144:16]
  assign io_fw_bottom_1 = fw_bottom_reg_1; // @[CrossBarSwitch.scala 144:16]
  assign io_fw_bottom_2 = fw_bottom_reg_2; // @[CrossBarSwitch.scala 144:16]
  assign io_fw_bottom_3 = fw_bottom_reg_3; // @[CrossBarSwitch.scala 144:16]
  assign cells_2d_0_io_fw_left = io_fw_left_0; // @[CrossBarSwitch.scala 126:29]
  assign cells_2d_0_io_fw_top = 65'h0; // @[CrossBarSwitch.scala 118:28]
  assign cells_2d_0_io_sel = select_onehot_0[0]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_1_io_fw_left = cells_2d_0_io_fw_right; // @[CrossBarSwitch.scala 129:29]
  assign cells_2d_1_io_fw_top = 65'h0; // @[CrossBarSwitch.scala 118:28]
  assign cells_2d_1_io_sel = select_onehot_1[0]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_2_io_fw_left = cells_2d_1_io_fw_right; // @[CrossBarSwitch.scala 129:29]
  assign cells_2d_2_io_fw_top = 65'h0; // @[CrossBarSwitch.scala 118:28]
  assign cells_2d_2_io_sel = select_onehot_2[0]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_3_io_fw_left = cells_2d_2_io_fw_right; // @[CrossBarSwitch.scala 129:29]
  assign cells_2d_3_io_fw_top = 65'h0; // @[CrossBarSwitch.scala 118:28]
  assign cells_2d_3_io_sel = select_onehot_3[0]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_4_io_fw_left = io_fw_left_1; // @[CrossBarSwitch.scala 126:29]
  assign cells_2d_4_io_fw_top = cells_2d_0_io_fw_bottom; // @[CrossBarSwitch.scala 121:28]
  assign cells_2d_4_io_sel = select_onehot_0[1]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_5_io_fw_left = cells_2d_4_io_fw_right; // @[CrossBarSwitch.scala 129:29]
  assign cells_2d_5_io_fw_top = cells_2d_1_io_fw_bottom; // @[CrossBarSwitch.scala 121:28]
  assign cells_2d_5_io_sel = select_onehot_1[1]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_6_io_fw_left = cells_2d_5_io_fw_right; // @[CrossBarSwitch.scala 129:29]
  assign cells_2d_6_io_fw_top = cells_2d_2_io_fw_bottom; // @[CrossBarSwitch.scala 121:28]
  assign cells_2d_6_io_sel = select_onehot_2[1]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_7_io_fw_left = cells_2d_6_io_fw_right; // @[CrossBarSwitch.scala 129:29]
  assign cells_2d_7_io_fw_top = cells_2d_3_io_fw_bottom; // @[CrossBarSwitch.scala 121:28]
  assign cells_2d_7_io_sel = select_onehot_3[1]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_8_io_fw_left = io_fw_left_2; // @[CrossBarSwitch.scala 126:29]
  assign cells_2d_8_io_fw_top = cells_2d_4_io_fw_bottom; // @[CrossBarSwitch.scala 121:28]
  assign cells_2d_8_io_sel = select_onehot_0[2]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_9_io_fw_left = cells_2d_8_io_fw_right; // @[CrossBarSwitch.scala 129:29]
  assign cells_2d_9_io_fw_top = cells_2d_5_io_fw_bottom; // @[CrossBarSwitch.scala 121:28]
  assign cells_2d_9_io_sel = select_onehot_1[2]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_10_io_fw_left = cells_2d_9_io_fw_right; // @[CrossBarSwitch.scala 129:29]
  assign cells_2d_10_io_fw_top = cells_2d_6_io_fw_bottom; // @[CrossBarSwitch.scala 121:28]
  assign cells_2d_10_io_sel = select_onehot_2[2]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_11_io_fw_left = cells_2d_10_io_fw_right; // @[CrossBarSwitch.scala 129:29]
  assign cells_2d_11_io_fw_top = cells_2d_7_io_fw_bottom; // @[CrossBarSwitch.scala 121:28]
  assign cells_2d_11_io_sel = select_onehot_3[2]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_12_io_fw_left = io_fw_left_3; // @[CrossBarSwitch.scala 126:29]
  assign cells_2d_12_io_fw_top = cells_2d_8_io_fw_bottom; // @[CrossBarSwitch.scala 121:28]
  assign cells_2d_12_io_sel = select_onehot_0[3]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_13_io_fw_left = cells_2d_12_io_fw_right; // @[CrossBarSwitch.scala 129:29]
  assign cells_2d_13_io_fw_top = cells_2d_9_io_fw_bottom; // @[CrossBarSwitch.scala 121:28]
  assign cells_2d_13_io_sel = select_onehot_1[3]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_14_io_fw_left = cells_2d_13_io_fw_right; // @[CrossBarSwitch.scala 129:29]
  assign cells_2d_14_io_fw_top = cells_2d_10_io_fw_bottom; // @[CrossBarSwitch.scala 121:28]
  assign cells_2d_14_io_sel = select_onehot_2[3]; // @[CrossBarSwitch.scala 133:44]
  assign cells_2d_15_io_fw_left = cells_2d_14_io_fw_right; // @[CrossBarSwitch.scala 129:29]
  assign cells_2d_15_io_fw_top = cells_2d_11_io_fw_bottom; // @[CrossBarSwitch.scala 121:28]
  assign cells_2d_15_io_sel = select_onehot_3[3]; // @[CrossBarSwitch.scala 133:44]
  always @(posedge clock) begin
    fw_bottom_reg_0 <= cells_2d_12_io_fw_bottom; // @[CrossBarSwitch.scala 141:22]
    fw_bottom_reg_1 <= cells_2d_13_io_fw_bottom; // @[CrossBarSwitch.scala 141:22]
    fw_bottom_reg_2 <= cells_2d_14_io_fw_bottom; // @[CrossBarSwitch.scala 141:22]
    fw_bottom_reg_3 <= cells_2d_15_io_fw_bottom; // @[CrossBarSwitch.scala 141:22]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  fw_bottom_reg_0 = _RAND_0[64:0];
  _RAND_1 = {3{`RANDOM}};
  fw_bottom_reg_1 = _RAND_1[64:0];
  _RAND_2 = {3{`RANDOM}};
  fw_bottom_reg_2 = _RAND_2[64:0];
  _RAND_3 = {3{`RANDOM}};
  fw_bottom_reg_3 = _RAND_3[64:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CLOScell4(
  input         clock,
  input  [64:0] io_in4_0,
  input  [64:0] io_in4_1,
  input  [64:0] io_in4_2,
  input  [64:0] io_in4_3,
  output [64:0] io_out4_0,
  output [64:0] io_out4_1,
  output [64:0] io_out4_2,
  output [64:0] io_out4_3,
  input  [7:0]  io_ctrl
);
  wire  CrossBarSwitch_clock; // @[BuildingBlock.scala 19:21]
  wire [64:0] CrossBarSwitch_io_fw_left_0; // @[BuildingBlock.scala 19:21]
  wire [64:0] CrossBarSwitch_io_fw_left_1; // @[BuildingBlock.scala 19:21]
  wire [64:0] CrossBarSwitch_io_fw_left_2; // @[BuildingBlock.scala 19:21]
  wire [64:0] CrossBarSwitch_io_fw_left_3; // @[BuildingBlock.scala 19:21]
  wire [64:0] CrossBarSwitch_io_fw_bottom_0; // @[BuildingBlock.scala 19:21]
  wire [64:0] CrossBarSwitch_io_fw_bottom_1; // @[BuildingBlock.scala 19:21]
  wire [64:0] CrossBarSwitch_io_fw_bottom_2; // @[BuildingBlock.scala 19:21]
  wire [64:0] CrossBarSwitch_io_fw_bottom_3; // @[BuildingBlock.scala 19:21]
  wire [1:0] CrossBarSwitch_io_select_0; // @[BuildingBlock.scala 19:21]
  wire [1:0] CrossBarSwitch_io_select_1; // @[BuildingBlock.scala 19:21]
  wire [1:0] CrossBarSwitch_io_select_2; // @[BuildingBlock.scala 19:21]
  wire [1:0] CrossBarSwitch_io_select_3; // @[BuildingBlock.scala 19:21]
  CrossBarSwitch CrossBarSwitch ( // @[BuildingBlock.scala 19:21]
    .clock(CrossBarSwitch_clock),
    .io_fw_left_0(CrossBarSwitch_io_fw_left_0),
    .io_fw_left_1(CrossBarSwitch_io_fw_left_1),
    .io_fw_left_2(CrossBarSwitch_io_fw_left_2),
    .io_fw_left_3(CrossBarSwitch_io_fw_left_3),
    .io_fw_bottom_0(CrossBarSwitch_io_fw_bottom_0),
    .io_fw_bottom_1(CrossBarSwitch_io_fw_bottom_1),
    .io_fw_bottom_2(CrossBarSwitch_io_fw_bottom_2),
    .io_fw_bottom_3(CrossBarSwitch_io_fw_bottom_3),
    .io_select_0(CrossBarSwitch_io_select_0),
    .io_select_1(CrossBarSwitch_io_select_1),
    .io_select_2(CrossBarSwitch_io_select_2),
    .io_select_3(CrossBarSwitch_io_select_3)
  );
  assign io_out4_0 = CrossBarSwitch_io_fw_bottom_0; // @[BuildingBlock.scala 24:11]
  assign io_out4_1 = CrossBarSwitch_io_fw_bottom_1; // @[BuildingBlock.scala 24:11]
  assign io_out4_2 = CrossBarSwitch_io_fw_bottom_2; // @[BuildingBlock.scala 24:11]
  assign io_out4_3 = CrossBarSwitch_io_fw_bottom_3; // @[BuildingBlock.scala 24:11]
  assign CrossBarSwitch_clock = clock;
  assign CrossBarSwitch_io_fw_left_0 = io_in4_0; // @[BuildingBlock.scala 23:17]
  assign CrossBarSwitch_io_fw_left_1 = io_in4_1; // @[BuildingBlock.scala 23:17]
  assign CrossBarSwitch_io_fw_left_2 = io_in4_2; // @[BuildingBlock.scala 23:17]
  assign CrossBarSwitch_io_fw_left_3 = io_in4_3; // @[BuildingBlock.scala 23:17]
  assign CrossBarSwitch_io_select_0 = io_ctrl[7:6]; // @[BuildingBlock.scala 21:31]
  assign CrossBarSwitch_io_select_1 = io_ctrl[5:4]; // @[BuildingBlock.scala 21:31]
  assign CrossBarSwitch_io_select_2 = io_ctrl[3:2]; // @[BuildingBlock.scala 21:31]
  assign CrossBarSwitch_io_select_3 = io_ctrl[1:0]; // @[BuildingBlock.scala 21:31]
endmodule
module CLOSingress1(
  input          clock,
  input  [63:0]  io_in64_0,
  input  [63:0]  io_in64_1,
  input  [63:0]  io_in64_2,
  input  [63:0]  io_in64_3,
  input  [63:0]  io_in64_4,
  input  [63:0]  io_in64_5,
  input  [63:0]  io_in64_6,
  input  [63:0]  io_in64_7,
  input  [63:0]  io_in64_8,
  input  [63:0]  io_in64_9,
  input  [63:0]  io_in64_10,
  input  [63:0]  io_in64_11,
  input  [63:0]  io_in64_12,
  input  [63:0]  io_in64_13,
  input  [63:0]  io_in64_14,
  input  [63:0]  io_in64_15,
  input  [63:0]  io_in64_16,
  input  [63:0]  io_in64_17,
  input  [63:0]  io_in64_18,
  input  [63:0]  io_in64_19,
  input  [63:0]  io_in64_20,
  input  [63:0]  io_in64_21,
  input  [63:0]  io_in64_22,
  input  [63:0]  io_in64_23,
  input  [63:0]  io_in64_24,
  input  [63:0]  io_in64_25,
  input  [63:0]  io_in64_26,
  input  [63:0]  io_in64_27,
  input  [63:0]  io_in64_28,
  input  [63:0]  io_in64_29,
  input  [63:0]  io_in64_30,
  input  [63:0]  io_in64_31,
  input  [63:0]  io_in64_32,
  input  [63:0]  io_in64_33,
  input  [63:0]  io_in64_34,
  input  [63:0]  io_in64_35,
  input  [63:0]  io_in64_36,
  input  [63:0]  io_in64_37,
  input  [63:0]  io_in64_38,
  input  [63:0]  io_in64_39,
  input  [63:0]  io_in64_40,
  input  [63:0]  io_in64_41,
  input  [63:0]  io_in64_42,
  input  [63:0]  io_in64_43,
  input  [63:0]  io_in64_44,
  input  [63:0]  io_in64_45,
  input  [63:0]  io_in64_46,
  input  [63:0]  io_in64_47,
  input  [63:0]  io_in64_48,
  input  [63:0]  io_in64_49,
  input  [63:0]  io_in64_50,
  input  [63:0]  io_in64_51,
  input  [63:0]  io_in64_52,
  input  [63:0]  io_in64_53,
  input  [63:0]  io_in64_54,
  input  [63:0]  io_in64_55,
  input  [63:0]  io_in64_56,
  input  [63:0]  io_in64_57,
  input  [63:0]  io_in64_58,
  input  [63:0]  io_in64_59,
  input  [63:0]  io_in64_60,
  input  [63:0]  io_in64_61,
  input  [63:0]  io_in64_62,
  input  [63:0]  io_in64_63,
  input          io_validin64_0,
  input          io_validin64_2,
  input          io_validin64_4,
  input          io_validin64_6,
  input          io_validin64_8,
  input          io_validin64_10,
  input          io_validin64_12,
  input          io_validin64_14,
  input          io_validin64_16,
  input          io_validin64_18,
  input          io_validin64_20,
  input          io_validin64_22,
  input          io_validin64_24,
  input          io_validin64_26,
  input          io_validin64_28,
  input          io_validin64_30,
  input          io_validin64_32,
  input          io_validin64_34,
  input          io_validin64_36,
  input          io_validin64_38,
  input          io_validin64_40,
  input          io_validin64_42,
  input          io_validin64_44,
  input          io_validin64_46,
  input          io_validin64_48,
  input          io_validin64_50,
  input          io_validin64_52,
  input          io_validin64_54,
  input          io_validin64_56,
  input          io_validin64_58,
  input          io_validin64_60,
  input          io_validin64_62,
  input  [1:0]   io_tagin_Tag,
  input  [2:0]   io_tagin_RoundCnt,
  input  [7:0]   io_addrin,
  output [63:0]  io_out64_0,
  output [63:0]  io_out64_1,
  output [63:0]  io_out64_2,
  output [63:0]  io_out64_3,
  output [63:0]  io_out64_4,
  output [63:0]  io_out64_5,
  output [63:0]  io_out64_6,
  output [63:0]  io_out64_7,
  output [63:0]  io_out64_8,
  output [63:0]  io_out64_9,
  output [63:0]  io_out64_10,
  output [63:0]  io_out64_11,
  output [63:0]  io_out64_12,
  output [63:0]  io_out64_13,
  output [63:0]  io_out64_14,
  output [63:0]  io_out64_15,
  output [63:0]  io_out64_16,
  output [63:0]  io_out64_17,
  output [63:0]  io_out64_18,
  output [63:0]  io_out64_19,
  output [63:0]  io_out64_20,
  output [63:0]  io_out64_21,
  output [63:0]  io_out64_22,
  output [63:0]  io_out64_23,
  output [63:0]  io_out64_24,
  output [63:0]  io_out64_25,
  output [63:0]  io_out64_26,
  output [63:0]  io_out64_27,
  output [63:0]  io_out64_28,
  output [63:0]  io_out64_29,
  output [63:0]  io_out64_30,
  output [63:0]  io_out64_31,
  output [63:0]  io_out64_32,
  output [63:0]  io_out64_33,
  output [63:0]  io_out64_34,
  output [63:0]  io_out64_35,
  output [63:0]  io_out64_36,
  output [63:0]  io_out64_37,
  output [63:0]  io_out64_38,
  output [63:0]  io_out64_39,
  output [63:0]  io_out64_40,
  output [63:0]  io_out64_41,
  output [63:0]  io_out64_42,
  output [63:0]  io_out64_43,
  output [63:0]  io_out64_44,
  output [63:0]  io_out64_45,
  output [63:0]  io_out64_46,
  output [63:0]  io_out64_47,
  output [63:0]  io_out64_48,
  output [63:0]  io_out64_49,
  output [63:0]  io_out64_50,
  output [63:0]  io_out64_51,
  output [63:0]  io_out64_52,
  output [63:0]  io_out64_53,
  output [63:0]  io_out64_54,
  output [63:0]  io_out64_55,
  output [63:0]  io_out64_56,
  output [63:0]  io_out64_57,
  output [63:0]  io_out64_58,
  output [63:0]  io_out64_59,
  output [63:0]  io_out64_60,
  output [63:0]  io_out64_61,
  output [63:0]  io_out64_62,
  output [63:0]  io_out64_63,
  output         io_validout64_0,
  output         io_validout64_1,
  output         io_validout64_2,
  output         io_validout64_3,
  output         io_validout64_4,
  output         io_validout64_5,
  output         io_validout64_6,
  output         io_validout64_7,
  output         io_validout64_8,
  output         io_validout64_9,
  output         io_validout64_10,
  output         io_validout64_11,
  output         io_validout64_12,
  output         io_validout64_13,
  output         io_validout64_14,
  output         io_validout64_15,
  output         io_validout64_16,
  output         io_validout64_17,
  output         io_validout64_18,
  output         io_validout64_19,
  output         io_validout64_20,
  output         io_validout64_21,
  output         io_validout64_22,
  output         io_validout64_23,
  output         io_validout64_24,
  output         io_validout64_25,
  output         io_validout64_26,
  output         io_validout64_27,
  output         io_validout64_28,
  output         io_validout64_29,
  output         io_validout64_30,
  output         io_validout64_31,
  output         io_validout64_32,
  output         io_validout64_33,
  output         io_validout64_34,
  output         io_validout64_35,
  output         io_validout64_36,
  output         io_validout64_37,
  output         io_validout64_38,
  output         io_validout64_39,
  output         io_validout64_40,
  output         io_validout64_41,
  output         io_validout64_42,
  output         io_validout64_43,
  output         io_validout64_44,
  output         io_validout64_45,
  output         io_validout64_46,
  output         io_validout64_47,
  output         io_validout64_48,
  output         io_validout64_49,
  output         io_validout64_50,
  output         io_validout64_51,
  output         io_validout64_52,
  output         io_validout64_53,
  output         io_validout64_54,
  output         io_validout64_55,
  output         io_validout64_56,
  output         io_validout64_57,
  output         io_validout64_58,
  output         io_validout64_59,
  output         io_validout64_60,
  output         io_validout64_61,
  output         io_validout64_62,
  output         io_validout64_63,
  output [1:0]   io_tagout_Tag,
  output [2:0]   io_tagout_RoundCnt,
  output [7:0]   io_addrout,
  input  [127:0] io_ctrl
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ingress1_0_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_0_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_0_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_0_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_0_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_0_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_0_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_0_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_0_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_0_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_1_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_1_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_1_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_1_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_1_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_1_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_1_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_1_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_1_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_1_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_2_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_2_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_2_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_2_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_2_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_2_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_2_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_2_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_2_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_2_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_3_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_3_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_3_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_3_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_3_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_3_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_3_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_3_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_3_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_3_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_4_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_4_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_4_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_4_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_4_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_4_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_4_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_4_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_4_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_4_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_5_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_5_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_5_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_5_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_5_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_5_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_5_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_5_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_5_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_5_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_6_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_6_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_6_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_6_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_6_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_6_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_6_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_6_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_6_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_6_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_7_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_7_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_7_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_7_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_7_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_7_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_7_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_7_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_7_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_7_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_8_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_8_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_8_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_8_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_8_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_8_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_8_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_8_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_8_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_8_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_9_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_9_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_9_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_9_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_9_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_9_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_9_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_9_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_9_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_9_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_10_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_10_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_10_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_10_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_10_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_10_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_10_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_10_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_10_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_10_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_11_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_11_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_11_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_11_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_11_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_11_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_11_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_11_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_11_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_11_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_12_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_12_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_12_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_12_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_12_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_12_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_12_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_12_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_12_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_12_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_13_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_13_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_13_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_13_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_13_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_13_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_13_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_13_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_13_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_13_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_14_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_14_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_14_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_14_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_14_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_14_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_14_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_14_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_14_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_14_io_ctrl; // @[BuildingBlock.scala 40:52]
  wire  ingress1_15_clock; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_15_io_in4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_15_io_in4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_15_io_in4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_15_io_in4_3; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_15_io_out4_0; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_15_io_out4_1; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_15_io_out4_2; // @[BuildingBlock.scala 40:52]
  wire [64:0] ingress1_15_io_out4_3; // @[BuildingBlock.scala 40:52]
  wire [7:0] ingress1_15_io_ctrl; // @[BuildingBlock.scala 40:52]
  reg [1:0] tag_Tag; // @[BuildingBlock.scala 41:20]
  reg [2:0] tag_RoundCnt; // @[BuildingBlock.scala 41:20]
  reg [7:0] addr; // @[BuildingBlock.scala 43:21]
  CLOScell4 ingress1_0 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_0_clock),
    .io_in4_0(ingress1_0_io_in4_0),
    .io_in4_1(ingress1_0_io_in4_1),
    .io_in4_2(ingress1_0_io_in4_2),
    .io_in4_3(ingress1_0_io_in4_3),
    .io_out4_0(ingress1_0_io_out4_0),
    .io_out4_1(ingress1_0_io_out4_1),
    .io_out4_2(ingress1_0_io_out4_2),
    .io_out4_3(ingress1_0_io_out4_3),
    .io_ctrl(ingress1_0_io_ctrl)
  );
  CLOScell4 ingress1_1 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_1_clock),
    .io_in4_0(ingress1_1_io_in4_0),
    .io_in4_1(ingress1_1_io_in4_1),
    .io_in4_2(ingress1_1_io_in4_2),
    .io_in4_3(ingress1_1_io_in4_3),
    .io_out4_0(ingress1_1_io_out4_0),
    .io_out4_1(ingress1_1_io_out4_1),
    .io_out4_2(ingress1_1_io_out4_2),
    .io_out4_3(ingress1_1_io_out4_3),
    .io_ctrl(ingress1_1_io_ctrl)
  );
  CLOScell4 ingress1_2 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_2_clock),
    .io_in4_0(ingress1_2_io_in4_0),
    .io_in4_1(ingress1_2_io_in4_1),
    .io_in4_2(ingress1_2_io_in4_2),
    .io_in4_3(ingress1_2_io_in4_3),
    .io_out4_0(ingress1_2_io_out4_0),
    .io_out4_1(ingress1_2_io_out4_1),
    .io_out4_2(ingress1_2_io_out4_2),
    .io_out4_3(ingress1_2_io_out4_3),
    .io_ctrl(ingress1_2_io_ctrl)
  );
  CLOScell4 ingress1_3 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_3_clock),
    .io_in4_0(ingress1_3_io_in4_0),
    .io_in4_1(ingress1_3_io_in4_1),
    .io_in4_2(ingress1_3_io_in4_2),
    .io_in4_3(ingress1_3_io_in4_3),
    .io_out4_0(ingress1_3_io_out4_0),
    .io_out4_1(ingress1_3_io_out4_1),
    .io_out4_2(ingress1_3_io_out4_2),
    .io_out4_3(ingress1_3_io_out4_3),
    .io_ctrl(ingress1_3_io_ctrl)
  );
  CLOScell4 ingress1_4 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_4_clock),
    .io_in4_0(ingress1_4_io_in4_0),
    .io_in4_1(ingress1_4_io_in4_1),
    .io_in4_2(ingress1_4_io_in4_2),
    .io_in4_3(ingress1_4_io_in4_3),
    .io_out4_0(ingress1_4_io_out4_0),
    .io_out4_1(ingress1_4_io_out4_1),
    .io_out4_2(ingress1_4_io_out4_2),
    .io_out4_3(ingress1_4_io_out4_3),
    .io_ctrl(ingress1_4_io_ctrl)
  );
  CLOScell4 ingress1_5 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_5_clock),
    .io_in4_0(ingress1_5_io_in4_0),
    .io_in4_1(ingress1_5_io_in4_1),
    .io_in4_2(ingress1_5_io_in4_2),
    .io_in4_3(ingress1_5_io_in4_3),
    .io_out4_0(ingress1_5_io_out4_0),
    .io_out4_1(ingress1_5_io_out4_1),
    .io_out4_2(ingress1_5_io_out4_2),
    .io_out4_3(ingress1_5_io_out4_3),
    .io_ctrl(ingress1_5_io_ctrl)
  );
  CLOScell4 ingress1_6 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_6_clock),
    .io_in4_0(ingress1_6_io_in4_0),
    .io_in4_1(ingress1_6_io_in4_1),
    .io_in4_2(ingress1_6_io_in4_2),
    .io_in4_3(ingress1_6_io_in4_3),
    .io_out4_0(ingress1_6_io_out4_0),
    .io_out4_1(ingress1_6_io_out4_1),
    .io_out4_2(ingress1_6_io_out4_2),
    .io_out4_3(ingress1_6_io_out4_3),
    .io_ctrl(ingress1_6_io_ctrl)
  );
  CLOScell4 ingress1_7 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_7_clock),
    .io_in4_0(ingress1_7_io_in4_0),
    .io_in4_1(ingress1_7_io_in4_1),
    .io_in4_2(ingress1_7_io_in4_2),
    .io_in4_3(ingress1_7_io_in4_3),
    .io_out4_0(ingress1_7_io_out4_0),
    .io_out4_1(ingress1_7_io_out4_1),
    .io_out4_2(ingress1_7_io_out4_2),
    .io_out4_3(ingress1_7_io_out4_3),
    .io_ctrl(ingress1_7_io_ctrl)
  );
  CLOScell4 ingress1_8 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_8_clock),
    .io_in4_0(ingress1_8_io_in4_0),
    .io_in4_1(ingress1_8_io_in4_1),
    .io_in4_2(ingress1_8_io_in4_2),
    .io_in4_3(ingress1_8_io_in4_3),
    .io_out4_0(ingress1_8_io_out4_0),
    .io_out4_1(ingress1_8_io_out4_1),
    .io_out4_2(ingress1_8_io_out4_2),
    .io_out4_3(ingress1_8_io_out4_3),
    .io_ctrl(ingress1_8_io_ctrl)
  );
  CLOScell4 ingress1_9 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_9_clock),
    .io_in4_0(ingress1_9_io_in4_0),
    .io_in4_1(ingress1_9_io_in4_1),
    .io_in4_2(ingress1_9_io_in4_2),
    .io_in4_3(ingress1_9_io_in4_3),
    .io_out4_0(ingress1_9_io_out4_0),
    .io_out4_1(ingress1_9_io_out4_1),
    .io_out4_2(ingress1_9_io_out4_2),
    .io_out4_3(ingress1_9_io_out4_3),
    .io_ctrl(ingress1_9_io_ctrl)
  );
  CLOScell4 ingress1_10 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_10_clock),
    .io_in4_0(ingress1_10_io_in4_0),
    .io_in4_1(ingress1_10_io_in4_1),
    .io_in4_2(ingress1_10_io_in4_2),
    .io_in4_3(ingress1_10_io_in4_3),
    .io_out4_0(ingress1_10_io_out4_0),
    .io_out4_1(ingress1_10_io_out4_1),
    .io_out4_2(ingress1_10_io_out4_2),
    .io_out4_3(ingress1_10_io_out4_3),
    .io_ctrl(ingress1_10_io_ctrl)
  );
  CLOScell4 ingress1_11 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_11_clock),
    .io_in4_0(ingress1_11_io_in4_0),
    .io_in4_1(ingress1_11_io_in4_1),
    .io_in4_2(ingress1_11_io_in4_2),
    .io_in4_3(ingress1_11_io_in4_3),
    .io_out4_0(ingress1_11_io_out4_0),
    .io_out4_1(ingress1_11_io_out4_1),
    .io_out4_2(ingress1_11_io_out4_2),
    .io_out4_3(ingress1_11_io_out4_3),
    .io_ctrl(ingress1_11_io_ctrl)
  );
  CLOScell4 ingress1_12 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_12_clock),
    .io_in4_0(ingress1_12_io_in4_0),
    .io_in4_1(ingress1_12_io_in4_1),
    .io_in4_2(ingress1_12_io_in4_2),
    .io_in4_3(ingress1_12_io_in4_3),
    .io_out4_0(ingress1_12_io_out4_0),
    .io_out4_1(ingress1_12_io_out4_1),
    .io_out4_2(ingress1_12_io_out4_2),
    .io_out4_3(ingress1_12_io_out4_3),
    .io_ctrl(ingress1_12_io_ctrl)
  );
  CLOScell4 ingress1_13 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_13_clock),
    .io_in4_0(ingress1_13_io_in4_0),
    .io_in4_1(ingress1_13_io_in4_1),
    .io_in4_2(ingress1_13_io_in4_2),
    .io_in4_3(ingress1_13_io_in4_3),
    .io_out4_0(ingress1_13_io_out4_0),
    .io_out4_1(ingress1_13_io_out4_1),
    .io_out4_2(ingress1_13_io_out4_2),
    .io_out4_3(ingress1_13_io_out4_3),
    .io_ctrl(ingress1_13_io_ctrl)
  );
  CLOScell4 ingress1_14 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_14_clock),
    .io_in4_0(ingress1_14_io_in4_0),
    .io_in4_1(ingress1_14_io_in4_1),
    .io_in4_2(ingress1_14_io_in4_2),
    .io_in4_3(ingress1_14_io_in4_3),
    .io_out4_0(ingress1_14_io_out4_0),
    .io_out4_1(ingress1_14_io_out4_1),
    .io_out4_2(ingress1_14_io_out4_2),
    .io_out4_3(ingress1_14_io_out4_3),
    .io_ctrl(ingress1_14_io_ctrl)
  );
  CLOScell4 ingress1_15 ( // @[BuildingBlock.scala 40:52]
    .clock(ingress1_15_clock),
    .io_in4_0(ingress1_15_io_in4_0),
    .io_in4_1(ingress1_15_io_in4_1),
    .io_in4_2(ingress1_15_io_in4_2),
    .io_in4_3(ingress1_15_io_in4_3),
    .io_out4_0(ingress1_15_io_out4_0),
    .io_out4_1(ingress1_15_io_out4_1),
    .io_out4_2(ingress1_15_io_out4_2),
    .io_out4_3(ingress1_15_io_out4_3),
    .io_ctrl(ingress1_15_io_ctrl)
  );
  assign io_out64_0 = ingress1_0_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_1 = ingress1_1_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_2 = ingress1_2_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_3 = ingress1_3_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_4 = ingress1_4_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_5 = ingress1_5_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_6 = ingress1_6_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_7 = ingress1_7_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_8 = ingress1_8_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_9 = ingress1_9_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_10 = ingress1_10_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_11 = ingress1_11_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_12 = ingress1_12_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_13 = ingress1_13_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_14 = ingress1_14_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_15 = ingress1_15_io_out4_0[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_16 = ingress1_0_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_17 = ingress1_1_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_18 = ingress1_2_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_19 = ingress1_3_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_20 = ingress1_4_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_21 = ingress1_5_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_22 = ingress1_6_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_23 = ingress1_7_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_24 = ingress1_8_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_25 = ingress1_9_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_26 = ingress1_10_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_27 = ingress1_11_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_28 = ingress1_12_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_29 = ingress1_13_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_30 = ingress1_14_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_31 = ingress1_15_io_out4_1[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_32 = ingress1_0_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_33 = ingress1_1_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_34 = ingress1_2_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_35 = ingress1_3_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_36 = ingress1_4_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_37 = ingress1_5_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_38 = ingress1_6_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_39 = ingress1_7_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_40 = ingress1_8_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_41 = ingress1_9_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_42 = ingress1_10_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_43 = ingress1_11_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_44 = ingress1_12_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_45 = ingress1_13_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_46 = ingress1_14_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_47 = ingress1_15_io_out4_2[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_48 = ingress1_0_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_49 = ingress1_1_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_50 = ingress1_2_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_51 = ingress1_3_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_52 = ingress1_4_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_53 = ingress1_5_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_54 = ingress1_6_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_55 = ingress1_7_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_56 = ingress1_8_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_57 = ingress1_9_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_58 = ingress1_10_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_59 = ingress1_11_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_60 = ingress1_12_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_61 = ingress1_13_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_62 = ingress1_14_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_out64_63 = ingress1_15_io_out4_3[63:0]; // @[BuildingBlock.scala 54:49]
  assign io_validout64_0 = ingress1_0_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_1 = ingress1_1_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_2 = ingress1_2_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_3 = ingress1_3_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_4 = ingress1_4_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_5 = ingress1_5_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_6 = ingress1_6_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_7 = ingress1_7_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_8 = ingress1_8_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_9 = ingress1_9_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_10 = ingress1_10_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_11 = ingress1_11_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_12 = ingress1_12_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_13 = ingress1_13_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_14 = ingress1_14_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_15 = ingress1_15_io_out4_0[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_16 = ingress1_0_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_17 = ingress1_1_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_18 = ingress1_2_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_19 = ingress1_3_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_20 = ingress1_4_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_21 = ingress1_5_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_22 = ingress1_6_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_23 = ingress1_7_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_24 = ingress1_8_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_25 = ingress1_9_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_26 = ingress1_10_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_27 = ingress1_11_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_28 = ingress1_12_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_29 = ingress1_13_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_30 = ingress1_14_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_31 = ingress1_15_io_out4_1[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_32 = ingress1_0_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_33 = ingress1_1_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_34 = ingress1_2_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_35 = ingress1_3_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_36 = ingress1_4_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_37 = ingress1_5_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_38 = ingress1_6_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_39 = ingress1_7_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_40 = ingress1_8_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_41 = ingress1_9_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_42 = ingress1_10_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_43 = ingress1_11_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_44 = ingress1_12_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_45 = ingress1_13_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_46 = ingress1_14_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_47 = ingress1_15_io_out4_2[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_48 = ingress1_0_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_49 = ingress1_1_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_50 = ingress1_2_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_51 = ingress1_3_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_52 = ingress1_4_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_53 = ingress1_5_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_54 = ingress1_6_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_55 = ingress1_7_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_56 = ingress1_8_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_57 = ingress1_9_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_58 = ingress1_10_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_59 = ingress1_11_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_60 = ingress1_12_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_61 = ingress1_13_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_62 = ingress1_14_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_validout64_63 = ingress1_15_io_out4_3[64]; // @[BuildingBlock.scala 55:54]
  assign io_tagout_Tag = tag_Tag; // @[BuildingBlock.scala 42:13]
  assign io_tagout_RoundCnt = tag_RoundCnt; // @[BuildingBlock.scala 42:13]
  assign io_addrout = addr; // @[BuildingBlock.scala 44:14]
  assign ingress1_0_clock = clock;
  assign ingress1_0_io_in4_0 = {io_validin64_0,io_in64_0}; // @[Cat.scala 30:58]
  assign ingress1_0_io_in4_1 = {1'h0,io_in64_1}; // @[Cat.scala 30:58]
  assign ingress1_0_io_in4_2 = {io_validin64_2,io_in64_2}; // @[Cat.scala 30:58]
  assign ingress1_0_io_in4_3 = {1'h0,io_in64_3}; // @[Cat.scala 30:58]
  assign ingress1_0_io_ctrl = io_ctrl[127:120]; // @[BuildingBlock.scala 59:35]
  assign ingress1_1_clock = clock;
  assign ingress1_1_io_in4_0 = {io_validin64_4,io_in64_4}; // @[Cat.scala 30:58]
  assign ingress1_1_io_in4_1 = {1'h0,io_in64_5}; // @[Cat.scala 30:58]
  assign ingress1_1_io_in4_2 = {io_validin64_6,io_in64_6}; // @[Cat.scala 30:58]
  assign ingress1_1_io_in4_3 = {1'h0,io_in64_7}; // @[Cat.scala 30:58]
  assign ingress1_1_io_ctrl = io_ctrl[119:112]; // @[BuildingBlock.scala 59:35]
  assign ingress1_2_clock = clock;
  assign ingress1_2_io_in4_0 = {io_validin64_8,io_in64_8}; // @[Cat.scala 30:58]
  assign ingress1_2_io_in4_1 = {1'h0,io_in64_9}; // @[Cat.scala 30:58]
  assign ingress1_2_io_in4_2 = {io_validin64_10,io_in64_10}; // @[Cat.scala 30:58]
  assign ingress1_2_io_in4_3 = {1'h0,io_in64_11}; // @[Cat.scala 30:58]
  assign ingress1_2_io_ctrl = io_ctrl[111:104]; // @[BuildingBlock.scala 59:35]
  assign ingress1_3_clock = clock;
  assign ingress1_3_io_in4_0 = {io_validin64_12,io_in64_12}; // @[Cat.scala 30:58]
  assign ingress1_3_io_in4_1 = {1'h0,io_in64_13}; // @[Cat.scala 30:58]
  assign ingress1_3_io_in4_2 = {io_validin64_14,io_in64_14}; // @[Cat.scala 30:58]
  assign ingress1_3_io_in4_3 = {1'h0,io_in64_15}; // @[Cat.scala 30:58]
  assign ingress1_3_io_ctrl = io_ctrl[103:96]; // @[BuildingBlock.scala 59:35]
  assign ingress1_4_clock = clock;
  assign ingress1_4_io_in4_0 = {io_validin64_16,io_in64_16}; // @[Cat.scala 30:58]
  assign ingress1_4_io_in4_1 = {1'h0,io_in64_17}; // @[Cat.scala 30:58]
  assign ingress1_4_io_in4_2 = {io_validin64_18,io_in64_18}; // @[Cat.scala 30:58]
  assign ingress1_4_io_in4_3 = {1'h0,io_in64_19}; // @[Cat.scala 30:58]
  assign ingress1_4_io_ctrl = io_ctrl[95:88]; // @[BuildingBlock.scala 59:35]
  assign ingress1_5_clock = clock;
  assign ingress1_5_io_in4_0 = {io_validin64_20,io_in64_20}; // @[Cat.scala 30:58]
  assign ingress1_5_io_in4_1 = {1'h0,io_in64_21}; // @[Cat.scala 30:58]
  assign ingress1_5_io_in4_2 = {io_validin64_22,io_in64_22}; // @[Cat.scala 30:58]
  assign ingress1_5_io_in4_3 = {1'h0,io_in64_23}; // @[Cat.scala 30:58]
  assign ingress1_5_io_ctrl = io_ctrl[87:80]; // @[BuildingBlock.scala 59:35]
  assign ingress1_6_clock = clock;
  assign ingress1_6_io_in4_0 = {io_validin64_24,io_in64_24}; // @[Cat.scala 30:58]
  assign ingress1_6_io_in4_1 = {1'h0,io_in64_25}; // @[Cat.scala 30:58]
  assign ingress1_6_io_in4_2 = {io_validin64_26,io_in64_26}; // @[Cat.scala 30:58]
  assign ingress1_6_io_in4_3 = {1'h0,io_in64_27}; // @[Cat.scala 30:58]
  assign ingress1_6_io_ctrl = io_ctrl[79:72]; // @[BuildingBlock.scala 59:35]
  assign ingress1_7_clock = clock;
  assign ingress1_7_io_in4_0 = {io_validin64_28,io_in64_28}; // @[Cat.scala 30:58]
  assign ingress1_7_io_in4_1 = {1'h0,io_in64_29}; // @[Cat.scala 30:58]
  assign ingress1_7_io_in4_2 = {io_validin64_30,io_in64_30}; // @[Cat.scala 30:58]
  assign ingress1_7_io_in4_3 = {1'h0,io_in64_31}; // @[Cat.scala 30:58]
  assign ingress1_7_io_ctrl = io_ctrl[71:64]; // @[BuildingBlock.scala 59:35]
  assign ingress1_8_clock = clock;
  assign ingress1_8_io_in4_0 = {io_validin64_32,io_in64_32}; // @[Cat.scala 30:58]
  assign ingress1_8_io_in4_1 = {1'h0,io_in64_33}; // @[Cat.scala 30:58]
  assign ingress1_8_io_in4_2 = {io_validin64_34,io_in64_34}; // @[Cat.scala 30:58]
  assign ingress1_8_io_in4_3 = {1'h0,io_in64_35}; // @[Cat.scala 30:58]
  assign ingress1_8_io_ctrl = io_ctrl[63:56]; // @[BuildingBlock.scala 59:35]
  assign ingress1_9_clock = clock;
  assign ingress1_9_io_in4_0 = {io_validin64_36,io_in64_36}; // @[Cat.scala 30:58]
  assign ingress1_9_io_in4_1 = {1'h0,io_in64_37}; // @[Cat.scala 30:58]
  assign ingress1_9_io_in4_2 = {io_validin64_38,io_in64_38}; // @[Cat.scala 30:58]
  assign ingress1_9_io_in4_3 = {1'h0,io_in64_39}; // @[Cat.scala 30:58]
  assign ingress1_9_io_ctrl = io_ctrl[55:48]; // @[BuildingBlock.scala 59:35]
  assign ingress1_10_clock = clock;
  assign ingress1_10_io_in4_0 = {io_validin64_40,io_in64_40}; // @[Cat.scala 30:58]
  assign ingress1_10_io_in4_1 = {1'h0,io_in64_41}; // @[Cat.scala 30:58]
  assign ingress1_10_io_in4_2 = {io_validin64_42,io_in64_42}; // @[Cat.scala 30:58]
  assign ingress1_10_io_in4_3 = {1'h0,io_in64_43}; // @[Cat.scala 30:58]
  assign ingress1_10_io_ctrl = io_ctrl[47:40]; // @[BuildingBlock.scala 59:35]
  assign ingress1_11_clock = clock;
  assign ingress1_11_io_in4_0 = {io_validin64_44,io_in64_44}; // @[Cat.scala 30:58]
  assign ingress1_11_io_in4_1 = {1'h0,io_in64_45}; // @[Cat.scala 30:58]
  assign ingress1_11_io_in4_2 = {io_validin64_46,io_in64_46}; // @[Cat.scala 30:58]
  assign ingress1_11_io_in4_3 = {1'h0,io_in64_47}; // @[Cat.scala 30:58]
  assign ingress1_11_io_ctrl = io_ctrl[39:32]; // @[BuildingBlock.scala 59:35]
  assign ingress1_12_clock = clock;
  assign ingress1_12_io_in4_0 = {io_validin64_48,io_in64_48}; // @[Cat.scala 30:58]
  assign ingress1_12_io_in4_1 = {1'h0,io_in64_49}; // @[Cat.scala 30:58]
  assign ingress1_12_io_in4_2 = {io_validin64_50,io_in64_50}; // @[Cat.scala 30:58]
  assign ingress1_12_io_in4_3 = {1'h0,io_in64_51}; // @[Cat.scala 30:58]
  assign ingress1_12_io_ctrl = io_ctrl[31:24]; // @[BuildingBlock.scala 59:35]
  assign ingress1_13_clock = clock;
  assign ingress1_13_io_in4_0 = {io_validin64_52,io_in64_52}; // @[Cat.scala 30:58]
  assign ingress1_13_io_in4_1 = {1'h0,io_in64_53}; // @[Cat.scala 30:58]
  assign ingress1_13_io_in4_2 = {io_validin64_54,io_in64_54}; // @[Cat.scala 30:58]
  assign ingress1_13_io_in4_3 = {1'h0,io_in64_55}; // @[Cat.scala 30:58]
  assign ingress1_13_io_ctrl = io_ctrl[23:16]; // @[BuildingBlock.scala 59:35]
  assign ingress1_14_clock = clock;
  assign ingress1_14_io_in4_0 = {io_validin64_56,io_in64_56}; // @[Cat.scala 30:58]
  assign ingress1_14_io_in4_1 = {1'h0,io_in64_57}; // @[Cat.scala 30:58]
  assign ingress1_14_io_in4_2 = {io_validin64_58,io_in64_58}; // @[Cat.scala 30:58]
  assign ingress1_14_io_in4_3 = {1'h0,io_in64_59}; // @[Cat.scala 30:58]
  assign ingress1_14_io_ctrl = io_ctrl[15:8]; // @[BuildingBlock.scala 59:35]
  assign ingress1_15_clock = clock;
  assign ingress1_15_io_in4_0 = {io_validin64_60,io_in64_60}; // @[Cat.scala 30:58]
  assign ingress1_15_io_in4_1 = {1'h0,io_in64_61}; // @[Cat.scala 30:58]
  assign ingress1_15_io_in4_2 = {io_validin64_62,io_in64_62}; // @[Cat.scala 30:58]
  assign ingress1_15_io_in4_3 = {1'h0,io_in64_63}; // @[Cat.scala 30:58]
  assign ingress1_15_io_ctrl = io_ctrl[7:0]; // @[BuildingBlock.scala 59:35]
  always @(posedge clock) begin
    tag_Tag <= io_tagin_Tag; // @[BuildingBlock.scala 41:20]
    tag_RoundCnt <= io_tagin_RoundCnt; // @[BuildingBlock.scala 41:20]
    addr <= io_addrin; // @[BuildingBlock.scala 43:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_Tag = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  tag_RoundCnt = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  addr = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CLOSingress2(
  input          clock,
  input  [63:0]  io_in64_0,
  input  [63:0]  io_in64_1,
  input  [63:0]  io_in64_2,
  input  [63:0]  io_in64_3,
  input  [63:0]  io_in64_4,
  input  [63:0]  io_in64_5,
  input  [63:0]  io_in64_6,
  input  [63:0]  io_in64_7,
  input  [63:0]  io_in64_8,
  input  [63:0]  io_in64_9,
  input  [63:0]  io_in64_10,
  input  [63:0]  io_in64_11,
  input  [63:0]  io_in64_12,
  input  [63:0]  io_in64_13,
  input  [63:0]  io_in64_14,
  input  [63:0]  io_in64_15,
  input  [63:0]  io_in64_16,
  input  [63:0]  io_in64_17,
  input  [63:0]  io_in64_18,
  input  [63:0]  io_in64_19,
  input  [63:0]  io_in64_20,
  input  [63:0]  io_in64_21,
  input  [63:0]  io_in64_22,
  input  [63:0]  io_in64_23,
  input  [63:0]  io_in64_24,
  input  [63:0]  io_in64_25,
  input  [63:0]  io_in64_26,
  input  [63:0]  io_in64_27,
  input  [63:0]  io_in64_28,
  input  [63:0]  io_in64_29,
  input  [63:0]  io_in64_30,
  input  [63:0]  io_in64_31,
  input  [63:0]  io_in64_32,
  input  [63:0]  io_in64_33,
  input  [63:0]  io_in64_34,
  input  [63:0]  io_in64_35,
  input  [63:0]  io_in64_36,
  input  [63:0]  io_in64_37,
  input  [63:0]  io_in64_38,
  input  [63:0]  io_in64_39,
  input  [63:0]  io_in64_40,
  input  [63:0]  io_in64_41,
  input  [63:0]  io_in64_42,
  input  [63:0]  io_in64_43,
  input  [63:0]  io_in64_44,
  input  [63:0]  io_in64_45,
  input  [63:0]  io_in64_46,
  input  [63:0]  io_in64_47,
  input  [63:0]  io_in64_48,
  input  [63:0]  io_in64_49,
  input  [63:0]  io_in64_50,
  input  [63:0]  io_in64_51,
  input  [63:0]  io_in64_52,
  input  [63:0]  io_in64_53,
  input  [63:0]  io_in64_54,
  input  [63:0]  io_in64_55,
  input  [63:0]  io_in64_56,
  input  [63:0]  io_in64_57,
  input  [63:0]  io_in64_58,
  input  [63:0]  io_in64_59,
  input  [63:0]  io_in64_60,
  input  [63:0]  io_in64_61,
  input  [63:0]  io_in64_62,
  input  [63:0]  io_in64_63,
  input          io_validin64_0,
  input          io_validin64_1,
  input          io_validin64_2,
  input          io_validin64_3,
  input          io_validin64_4,
  input          io_validin64_5,
  input          io_validin64_6,
  input          io_validin64_7,
  input          io_validin64_8,
  input          io_validin64_9,
  input          io_validin64_10,
  input          io_validin64_11,
  input          io_validin64_12,
  input          io_validin64_13,
  input          io_validin64_14,
  input          io_validin64_15,
  input          io_validin64_16,
  input          io_validin64_17,
  input          io_validin64_18,
  input          io_validin64_19,
  input          io_validin64_20,
  input          io_validin64_21,
  input          io_validin64_22,
  input          io_validin64_23,
  input          io_validin64_24,
  input          io_validin64_25,
  input          io_validin64_26,
  input          io_validin64_27,
  input          io_validin64_28,
  input          io_validin64_29,
  input          io_validin64_30,
  input          io_validin64_31,
  input          io_validin64_32,
  input          io_validin64_33,
  input          io_validin64_34,
  input          io_validin64_35,
  input          io_validin64_36,
  input          io_validin64_37,
  input          io_validin64_38,
  input          io_validin64_39,
  input          io_validin64_40,
  input          io_validin64_41,
  input          io_validin64_42,
  input          io_validin64_43,
  input          io_validin64_44,
  input          io_validin64_45,
  input          io_validin64_46,
  input          io_validin64_47,
  input          io_validin64_48,
  input          io_validin64_49,
  input          io_validin64_50,
  input          io_validin64_51,
  input          io_validin64_52,
  input          io_validin64_53,
  input          io_validin64_54,
  input          io_validin64_55,
  input          io_validin64_56,
  input          io_validin64_57,
  input          io_validin64_58,
  input          io_validin64_59,
  input          io_validin64_60,
  input          io_validin64_61,
  input          io_validin64_62,
  input          io_validin64_63,
  input  [1:0]   io_tagin_Tag,
  input  [2:0]   io_tagin_RoundCnt,
  input  [7:0]   io_addrin,
  output [63:0]  io_out64_0,
  output [63:0]  io_out64_1,
  output [63:0]  io_out64_2,
  output [63:0]  io_out64_3,
  output [63:0]  io_out64_4,
  output [63:0]  io_out64_5,
  output [63:0]  io_out64_6,
  output [63:0]  io_out64_7,
  output [63:0]  io_out64_8,
  output [63:0]  io_out64_9,
  output [63:0]  io_out64_10,
  output [63:0]  io_out64_11,
  output [63:0]  io_out64_12,
  output [63:0]  io_out64_13,
  output [63:0]  io_out64_14,
  output [63:0]  io_out64_15,
  output [63:0]  io_out64_16,
  output [63:0]  io_out64_17,
  output [63:0]  io_out64_18,
  output [63:0]  io_out64_19,
  output [63:0]  io_out64_20,
  output [63:0]  io_out64_21,
  output [63:0]  io_out64_22,
  output [63:0]  io_out64_23,
  output [63:0]  io_out64_24,
  output [63:0]  io_out64_25,
  output [63:0]  io_out64_26,
  output [63:0]  io_out64_27,
  output [63:0]  io_out64_28,
  output [63:0]  io_out64_29,
  output [63:0]  io_out64_30,
  output [63:0]  io_out64_31,
  output [63:0]  io_out64_32,
  output [63:0]  io_out64_33,
  output [63:0]  io_out64_34,
  output [63:0]  io_out64_35,
  output [63:0]  io_out64_36,
  output [63:0]  io_out64_37,
  output [63:0]  io_out64_38,
  output [63:0]  io_out64_39,
  output [63:0]  io_out64_40,
  output [63:0]  io_out64_41,
  output [63:0]  io_out64_42,
  output [63:0]  io_out64_43,
  output [63:0]  io_out64_44,
  output [63:0]  io_out64_45,
  output [63:0]  io_out64_46,
  output [63:0]  io_out64_47,
  output [63:0]  io_out64_48,
  output [63:0]  io_out64_49,
  output [63:0]  io_out64_50,
  output [63:0]  io_out64_51,
  output [63:0]  io_out64_52,
  output [63:0]  io_out64_53,
  output [63:0]  io_out64_54,
  output [63:0]  io_out64_55,
  output [63:0]  io_out64_56,
  output [63:0]  io_out64_57,
  output [63:0]  io_out64_58,
  output [63:0]  io_out64_59,
  output [63:0]  io_out64_60,
  output [63:0]  io_out64_61,
  output [63:0]  io_out64_62,
  output [63:0]  io_out64_63,
  output         io_validout64_0,
  output         io_validout64_1,
  output         io_validout64_2,
  output         io_validout64_3,
  output         io_validout64_4,
  output         io_validout64_5,
  output         io_validout64_6,
  output         io_validout64_7,
  output         io_validout64_8,
  output         io_validout64_9,
  output         io_validout64_10,
  output         io_validout64_11,
  output         io_validout64_12,
  output         io_validout64_13,
  output         io_validout64_14,
  output         io_validout64_15,
  output         io_validout64_16,
  output         io_validout64_17,
  output         io_validout64_18,
  output         io_validout64_19,
  output         io_validout64_20,
  output         io_validout64_21,
  output         io_validout64_22,
  output         io_validout64_23,
  output         io_validout64_24,
  output         io_validout64_25,
  output         io_validout64_26,
  output         io_validout64_27,
  output         io_validout64_28,
  output         io_validout64_29,
  output         io_validout64_30,
  output         io_validout64_31,
  output         io_validout64_32,
  output         io_validout64_33,
  output         io_validout64_34,
  output         io_validout64_35,
  output         io_validout64_36,
  output         io_validout64_37,
  output         io_validout64_38,
  output         io_validout64_39,
  output         io_validout64_40,
  output         io_validout64_41,
  output         io_validout64_42,
  output         io_validout64_43,
  output         io_validout64_44,
  output         io_validout64_45,
  output         io_validout64_46,
  output         io_validout64_47,
  output         io_validout64_48,
  output         io_validout64_49,
  output         io_validout64_50,
  output         io_validout64_51,
  output         io_validout64_52,
  output         io_validout64_53,
  output         io_validout64_54,
  output         io_validout64_55,
  output         io_validout64_56,
  output         io_validout64_57,
  output         io_validout64_58,
  output         io_validout64_59,
  output         io_validout64_60,
  output         io_validout64_61,
  output         io_validout64_62,
  output         io_validout64_63,
  output [1:0]   io_tagout_Tag,
  output [2:0]   io_tagout_RoundCnt,
  output [7:0]   io_addrout,
  input  [127:0] io_ctrl
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  ingress2_0_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_0_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_0_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_0_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_0_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_0_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_0_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_0_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_0_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_0_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_1_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_1_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_1_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_1_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_1_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_1_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_1_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_1_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_1_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_1_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_2_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_2_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_2_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_2_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_2_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_2_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_2_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_2_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_2_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_2_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_3_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_3_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_3_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_3_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_3_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_3_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_3_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_3_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_3_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_3_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_4_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_4_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_4_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_4_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_4_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_4_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_4_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_4_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_4_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_4_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_5_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_5_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_5_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_5_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_5_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_5_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_5_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_5_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_5_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_5_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_6_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_6_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_6_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_6_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_6_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_6_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_6_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_6_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_6_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_6_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_7_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_7_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_7_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_7_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_7_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_7_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_7_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_7_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_7_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_7_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_8_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_8_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_8_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_8_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_8_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_8_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_8_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_8_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_8_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_8_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_9_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_9_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_9_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_9_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_9_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_9_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_9_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_9_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_9_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_9_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_10_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_10_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_10_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_10_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_10_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_10_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_10_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_10_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_10_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_10_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_11_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_11_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_11_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_11_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_11_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_11_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_11_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_11_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_11_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_11_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_12_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_12_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_12_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_12_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_12_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_12_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_12_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_12_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_12_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_12_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_13_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_13_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_13_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_13_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_13_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_13_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_13_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_13_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_13_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_13_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_14_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_14_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_14_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_14_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_14_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_14_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_14_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_14_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_14_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_14_io_ctrl; // @[BuildingBlock.scala 75:52]
  wire  ingress2_15_clock; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_15_io_in4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_15_io_in4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_15_io_in4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_15_io_in4_3; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_15_io_out4_0; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_15_io_out4_1; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_15_io_out4_2; // @[BuildingBlock.scala 75:52]
  wire [64:0] ingress2_15_io_out4_3; // @[BuildingBlock.scala 75:52]
  wire [7:0] ingress2_15_io_ctrl; // @[BuildingBlock.scala 75:52]
  reg [1:0] tag_Tag; // @[BuildingBlock.scala 76:20]
  reg [2:0] tag_RoundCnt; // @[BuildingBlock.scala 76:20]
  reg [7:0] addr; // @[BuildingBlock.scala 78:21]
  CLOScell4 ingress2_0 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_0_clock),
    .io_in4_0(ingress2_0_io_in4_0),
    .io_in4_1(ingress2_0_io_in4_1),
    .io_in4_2(ingress2_0_io_in4_2),
    .io_in4_3(ingress2_0_io_in4_3),
    .io_out4_0(ingress2_0_io_out4_0),
    .io_out4_1(ingress2_0_io_out4_1),
    .io_out4_2(ingress2_0_io_out4_2),
    .io_out4_3(ingress2_0_io_out4_3),
    .io_ctrl(ingress2_0_io_ctrl)
  );
  CLOScell4 ingress2_1 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_1_clock),
    .io_in4_0(ingress2_1_io_in4_0),
    .io_in4_1(ingress2_1_io_in4_1),
    .io_in4_2(ingress2_1_io_in4_2),
    .io_in4_3(ingress2_1_io_in4_3),
    .io_out4_0(ingress2_1_io_out4_0),
    .io_out4_1(ingress2_1_io_out4_1),
    .io_out4_2(ingress2_1_io_out4_2),
    .io_out4_3(ingress2_1_io_out4_3),
    .io_ctrl(ingress2_1_io_ctrl)
  );
  CLOScell4 ingress2_2 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_2_clock),
    .io_in4_0(ingress2_2_io_in4_0),
    .io_in4_1(ingress2_2_io_in4_1),
    .io_in4_2(ingress2_2_io_in4_2),
    .io_in4_3(ingress2_2_io_in4_3),
    .io_out4_0(ingress2_2_io_out4_0),
    .io_out4_1(ingress2_2_io_out4_1),
    .io_out4_2(ingress2_2_io_out4_2),
    .io_out4_3(ingress2_2_io_out4_3),
    .io_ctrl(ingress2_2_io_ctrl)
  );
  CLOScell4 ingress2_3 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_3_clock),
    .io_in4_0(ingress2_3_io_in4_0),
    .io_in4_1(ingress2_3_io_in4_1),
    .io_in4_2(ingress2_3_io_in4_2),
    .io_in4_3(ingress2_3_io_in4_3),
    .io_out4_0(ingress2_3_io_out4_0),
    .io_out4_1(ingress2_3_io_out4_1),
    .io_out4_2(ingress2_3_io_out4_2),
    .io_out4_3(ingress2_3_io_out4_3),
    .io_ctrl(ingress2_3_io_ctrl)
  );
  CLOScell4 ingress2_4 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_4_clock),
    .io_in4_0(ingress2_4_io_in4_0),
    .io_in4_1(ingress2_4_io_in4_1),
    .io_in4_2(ingress2_4_io_in4_2),
    .io_in4_3(ingress2_4_io_in4_3),
    .io_out4_0(ingress2_4_io_out4_0),
    .io_out4_1(ingress2_4_io_out4_1),
    .io_out4_2(ingress2_4_io_out4_2),
    .io_out4_3(ingress2_4_io_out4_3),
    .io_ctrl(ingress2_4_io_ctrl)
  );
  CLOScell4 ingress2_5 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_5_clock),
    .io_in4_0(ingress2_5_io_in4_0),
    .io_in4_1(ingress2_5_io_in4_1),
    .io_in4_2(ingress2_5_io_in4_2),
    .io_in4_3(ingress2_5_io_in4_3),
    .io_out4_0(ingress2_5_io_out4_0),
    .io_out4_1(ingress2_5_io_out4_1),
    .io_out4_2(ingress2_5_io_out4_2),
    .io_out4_3(ingress2_5_io_out4_3),
    .io_ctrl(ingress2_5_io_ctrl)
  );
  CLOScell4 ingress2_6 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_6_clock),
    .io_in4_0(ingress2_6_io_in4_0),
    .io_in4_1(ingress2_6_io_in4_1),
    .io_in4_2(ingress2_6_io_in4_2),
    .io_in4_3(ingress2_6_io_in4_3),
    .io_out4_0(ingress2_6_io_out4_0),
    .io_out4_1(ingress2_6_io_out4_1),
    .io_out4_2(ingress2_6_io_out4_2),
    .io_out4_3(ingress2_6_io_out4_3),
    .io_ctrl(ingress2_6_io_ctrl)
  );
  CLOScell4 ingress2_7 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_7_clock),
    .io_in4_0(ingress2_7_io_in4_0),
    .io_in4_1(ingress2_7_io_in4_1),
    .io_in4_2(ingress2_7_io_in4_2),
    .io_in4_3(ingress2_7_io_in4_3),
    .io_out4_0(ingress2_7_io_out4_0),
    .io_out4_1(ingress2_7_io_out4_1),
    .io_out4_2(ingress2_7_io_out4_2),
    .io_out4_3(ingress2_7_io_out4_3),
    .io_ctrl(ingress2_7_io_ctrl)
  );
  CLOScell4 ingress2_8 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_8_clock),
    .io_in4_0(ingress2_8_io_in4_0),
    .io_in4_1(ingress2_8_io_in4_1),
    .io_in4_2(ingress2_8_io_in4_2),
    .io_in4_3(ingress2_8_io_in4_3),
    .io_out4_0(ingress2_8_io_out4_0),
    .io_out4_1(ingress2_8_io_out4_1),
    .io_out4_2(ingress2_8_io_out4_2),
    .io_out4_3(ingress2_8_io_out4_3),
    .io_ctrl(ingress2_8_io_ctrl)
  );
  CLOScell4 ingress2_9 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_9_clock),
    .io_in4_0(ingress2_9_io_in4_0),
    .io_in4_1(ingress2_9_io_in4_1),
    .io_in4_2(ingress2_9_io_in4_2),
    .io_in4_3(ingress2_9_io_in4_3),
    .io_out4_0(ingress2_9_io_out4_0),
    .io_out4_1(ingress2_9_io_out4_1),
    .io_out4_2(ingress2_9_io_out4_2),
    .io_out4_3(ingress2_9_io_out4_3),
    .io_ctrl(ingress2_9_io_ctrl)
  );
  CLOScell4 ingress2_10 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_10_clock),
    .io_in4_0(ingress2_10_io_in4_0),
    .io_in4_1(ingress2_10_io_in4_1),
    .io_in4_2(ingress2_10_io_in4_2),
    .io_in4_3(ingress2_10_io_in4_3),
    .io_out4_0(ingress2_10_io_out4_0),
    .io_out4_1(ingress2_10_io_out4_1),
    .io_out4_2(ingress2_10_io_out4_2),
    .io_out4_3(ingress2_10_io_out4_3),
    .io_ctrl(ingress2_10_io_ctrl)
  );
  CLOScell4 ingress2_11 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_11_clock),
    .io_in4_0(ingress2_11_io_in4_0),
    .io_in4_1(ingress2_11_io_in4_1),
    .io_in4_2(ingress2_11_io_in4_2),
    .io_in4_3(ingress2_11_io_in4_3),
    .io_out4_0(ingress2_11_io_out4_0),
    .io_out4_1(ingress2_11_io_out4_1),
    .io_out4_2(ingress2_11_io_out4_2),
    .io_out4_3(ingress2_11_io_out4_3),
    .io_ctrl(ingress2_11_io_ctrl)
  );
  CLOScell4 ingress2_12 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_12_clock),
    .io_in4_0(ingress2_12_io_in4_0),
    .io_in4_1(ingress2_12_io_in4_1),
    .io_in4_2(ingress2_12_io_in4_2),
    .io_in4_3(ingress2_12_io_in4_3),
    .io_out4_0(ingress2_12_io_out4_0),
    .io_out4_1(ingress2_12_io_out4_1),
    .io_out4_2(ingress2_12_io_out4_2),
    .io_out4_3(ingress2_12_io_out4_3),
    .io_ctrl(ingress2_12_io_ctrl)
  );
  CLOScell4 ingress2_13 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_13_clock),
    .io_in4_0(ingress2_13_io_in4_0),
    .io_in4_1(ingress2_13_io_in4_1),
    .io_in4_2(ingress2_13_io_in4_2),
    .io_in4_3(ingress2_13_io_in4_3),
    .io_out4_0(ingress2_13_io_out4_0),
    .io_out4_1(ingress2_13_io_out4_1),
    .io_out4_2(ingress2_13_io_out4_2),
    .io_out4_3(ingress2_13_io_out4_3),
    .io_ctrl(ingress2_13_io_ctrl)
  );
  CLOScell4 ingress2_14 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_14_clock),
    .io_in4_0(ingress2_14_io_in4_0),
    .io_in4_1(ingress2_14_io_in4_1),
    .io_in4_2(ingress2_14_io_in4_2),
    .io_in4_3(ingress2_14_io_in4_3),
    .io_out4_0(ingress2_14_io_out4_0),
    .io_out4_1(ingress2_14_io_out4_1),
    .io_out4_2(ingress2_14_io_out4_2),
    .io_out4_3(ingress2_14_io_out4_3),
    .io_ctrl(ingress2_14_io_ctrl)
  );
  CLOScell4 ingress2_15 ( // @[BuildingBlock.scala 75:52]
    .clock(ingress2_15_clock),
    .io_in4_0(ingress2_15_io_in4_0),
    .io_in4_1(ingress2_15_io_in4_1),
    .io_in4_2(ingress2_15_io_in4_2),
    .io_in4_3(ingress2_15_io_in4_3),
    .io_out4_0(ingress2_15_io_out4_0),
    .io_out4_1(ingress2_15_io_out4_1),
    .io_out4_2(ingress2_15_io_out4_2),
    .io_out4_3(ingress2_15_io_out4_3),
    .io_ctrl(ingress2_15_io_ctrl)
  );
  assign io_out64_0 = ingress2_0_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_1 = ingress2_1_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_2 = ingress2_2_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_3 = ingress2_3_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_4 = ingress2_0_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_5 = ingress2_1_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_6 = ingress2_2_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_7 = ingress2_3_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_8 = ingress2_0_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_9 = ingress2_1_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_10 = ingress2_2_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_11 = ingress2_3_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_12 = ingress2_0_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_13 = ingress2_1_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_14 = ingress2_2_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_15 = ingress2_3_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_16 = ingress2_4_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_17 = ingress2_5_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_18 = ingress2_6_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_19 = ingress2_7_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_20 = ingress2_4_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_21 = ingress2_5_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_22 = ingress2_6_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_23 = ingress2_7_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_24 = ingress2_4_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_25 = ingress2_5_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_26 = ingress2_6_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_27 = ingress2_7_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_28 = ingress2_4_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_29 = ingress2_5_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_30 = ingress2_6_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_31 = ingress2_7_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_32 = ingress2_8_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_33 = ingress2_9_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_34 = ingress2_10_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_35 = ingress2_11_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_36 = ingress2_8_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_37 = ingress2_9_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_38 = ingress2_10_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_39 = ingress2_11_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_40 = ingress2_8_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_41 = ingress2_9_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_42 = ingress2_10_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_43 = ingress2_11_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_44 = ingress2_8_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_45 = ingress2_9_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_46 = ingress2_10_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_47 = ingress2_11_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_48 = ingress2_12_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_49 = ingress2_13_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_50 = ingress2_14_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_51 = ingress2_15_io_out4_0[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_52 = ingress2_12_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_53 = ingress2_13_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_54 = ingress2_14_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_55 = ingress2_15_io_out4_1[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_56 = ingress2_12_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_57 = ingress2_13_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_58 = ingress2_14_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_59 = ingress2_15_io_out4_2[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_60 = ingress2_12_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_61 = ingress2_13_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_62 = ingress2_14_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_out64_63 = ingress2_15_io_out4_3[63:0]; // @[BuildingBlock.scala 90:59]
  assign io_validout64_0 = ingress2_0_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_1 = ingress2_1_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_2 = ingress2_2_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_3 = ingress2_3_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_4 = ingress2_0_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_5 = ingress2_1_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_6 = ingress2_2_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_7 = ingress2_3_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_8 = ingress2_0_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_9 = ingress2_1_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_10 = ingress2_2_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_11 = ingress2_3_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_12 = ingress2_0_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_13 = ingress2_1_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_14 = ingress2_2_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_15 = ingress2_3_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_16 = ingress2_4_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_17 = ingress2_5_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_18 = ingress2_6_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_19 = ingress2_7_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_20 = ingress2_4_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_21 = ingress2_5_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_22 = ingress2_6_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_23 = ingress2_7_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_24 = ingress2_4_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_25 = ingress2_5_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_26 = ingress2_6_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_27 = ingress2_7_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_28 = ingress2_4_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_29 = ingress2_5_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_30 = ingress2_6_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_31 = ingress2_7_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_32 = ingress2_8_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_33 = ingress2_9_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_34 = ingress2_10_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_35 = ingress2_11_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_36 = ingress2_8_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_37 = ingress2_9_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_38 = ingress2_10_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_39 = ingress2_11_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_40 = ingress2_8_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_41 = ingress2_9_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_42 = ingress2_10_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_43 = ingress2_11_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_44 = ingress2_8_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_45 = ingress2_9_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_46 = ingress2_10_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_47 = ingress2_11_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_48 = ingress2_12_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_49 = ingress2_13_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_50 = ingress2_14_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_51 = ingress2_15_io_out4_0[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_52 = ingress2_12_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_53 = ingress2_13_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_54 = ingress2_14_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_55 = ingress2_15_io_out4_1[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_56 = ingress2_12_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_57 = ingress2_13_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_58 = ingress2_14_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_59 = ingress2_15_io_out4_2[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_60 = ingress2_12_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_61 = ingress2_13_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_62 = ingress2_14_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_validout64_63 = ingress2_15_io_out4_3[64]; // @[BuildingBlock.scala 91:64]
  assign io_tagout_Tag = tag_Tag; // @[BuildingBlock.scala 77:13]
  assign io_tagout_RoundCnt = tag_RoundCnt; // @[BuildingBlock.scala 77:13]
  assign io_addrout = addr; // @[BuildingBlock.scala 79:14]
  assign ingress2_0_clock = clock;
  assign ingress2_0_io_in4_0 = {io_validin64_0,io_in64_0}; // @[Cat.scala 30:58]
  assign ingress2_0_io_in4_1 = {io_validin64_1,io_in64_1}; // @[Cat.scala 30:58]
  assign ingress2_0_io_in4_2 = {io_validin64_2,io_in64_2}; // @[Cat.scala 30:58]
  assign ingress2_0_io_in4_3 = {io_validin64_3,io_in64_3}; // @[Cat.scala 30:58]
  assign ingress2_0_io_ctrl = io_ctrl[127:120]; // @[BuildingBlock.scala 95:35]
  assign ingress2_1_clock = clock;
  assign ingress2_1_io_in4_0 = {io_validin64_4,io_in64_4}; // @[Cat.scala 30:58]
  assign ingress2_1_io_in4_1 = {io_validin64_5,io_in64_5}; // @[Cat.scala 30:58]
  assign ingress2_1_io_in4_2 = {io_validin64_6,io_in64_6}; // @[Cat.scala 30:58]
  assign ingress2_1_io_in4_3 = {io_validin64_7,io_in64_7}; // @[Cat.scala 30:58]
  assign ingress2_1_io_ctrl = io_ctrl[119:112]; // @[BuildingBlock.scala 95:35]
  assign ingress2_2_clock = clock;
  assign ingress2_2_io_in4_0 = {io_validin64_8,io_in64_8}; // @[Cat.scala 30:58]
  assign ingress2_2_io_in4_1 = {io_validin64_9,io_in64_9}; // @[Cat.scala 30:58]
  assign ingress2_2_io_in4_2 = {io_validin64_10,io_in64_10}; // @[Cat.scala 30:58]
  assign ingress2_2_io_in4_3 = {io_validin64_11,io_in64_11}; // @[Cat.scala 30:58]
  assign ingress2_2_io_ctrl = io_ctrl[111:104]; // @[BuildingBlock.scala 95:35]
  assign ingress2_3_clock = clock;
  assign ingress2_3_io_in4_0 = {io_validin64_12,io_in64_12}; // @[Cat.scala 30:58]
  assign ingress2_3_io_in4_1 = {io_validin64_13,io_in64_13}; // @[Cat.scala 30:58]
  assign ingress2_3_io_in4_2 = {io_validin64_14,io_in64_14}; // @[Cat.scala 30:58]
  assign ingress2_3_io_in4_3 = {io_validin64_15,io_in64_15}; // @[Cat.scala 30:58]
  assign ingress2_3_io_ctrl = io_ctrl[103:96]; // @[BuildingBlock.scala 95:35]
  assign ingress2_4_clock = clock;
  assign ingress2_4_io_in4_0 = {io_validin64_16,io_in64_16}; // @[Cat.scala 30:58]
  assign ingress2_4_io_in4_1 = {io_validin64_17,io_in64_17}; // @[Cat.scala 30:58]
  assign ingress2_4_io_in4_2 = {io_validin64_18,io_in64_18}; // @[Cat.scala 30:58]
  assign ingress2_4_io_in4_3 = {io_validin64_19,io_in64_19}; // @[Cat.scala 30:58]
  assign ingress2_4_io_ctrl = io_ctrl[95:88]; // @[BuildingBlock.scala 95:35]
  assign ingress2_5_clock = clock;
  assign ingress2_5_io_in4_0 = {io_validin64_20,io_in64_20}; // @[Cat.scala 30:58]
  assign ingress2_5_io_in4_1 = {io_validin64_21,io_in64_21}; // @[Cat.scala 30:58]
  assign ingress2_5_io_in4_2 = {io_validin64_22,io_in64_22}; // @[Cat.scala 30:58]
  assign ingress2_5_io_in4_3 = {io_validin64_23,io_in64_23}; // @[Cat.scala 30:58]
  assign ingress2_5_io_ctrl = io_ctrl[87:80]; // @[BuildingBlock.scala 95:35]
  assign ingress2_6_clock = clock;
  assign ingress2_6_io_in4_0 = {io_validin64_24,io_in64_24}; // @[Cat.scala 30:58]
  assign ingress2_6_io_in4_1 = {io_validin64_25,io_in64_25}; // @[Cat.scala 30:58]
  assign ingress2_6_io_in4_2 = {io_validin64_26,io_in64_26}; // @[Cat.scala 30:58]
  assign ingress2_6_io_in4_3 = {io_validin64_27,io_in64_27}; // @[Cat.scala 30:58]
  assign ingress2_6_io_ctrl = io_ctrl[79:72]; // @[BuildingBlock.scala 95:35]
  assign ingress2_7_clock = clock;
  assign ingress2_7_io_in4_0 = {io_validin64_28,io_in64_28}; // @[Cat.scala 30:58]
  assign ingress2_7_io_in4_1 = {io_validin64_29,io_in64_29}; // @[Cat.scala 30:58]
  assign ingress2_7_io_in4_2 = {io_validin64_30,io_in64_30}; // @[Cat.scala 30:58]
  assign ingress2_7_io_in4_3 = {io_validin64_31,io_in64_31}; // @[Cat.scala 30:58]
  assign ingress2_7_io_ctrl = io_ctrl[71:64]; // @[BuildingBlock.scala 95:35]
  assign ingress2_8_clock = clock;
  assign ingress2_8_io_in4_0 = {io_validin64_32,io_in64_32}; // @[Cat.scala 30:58]
  assign ingress2_8_io_in4_1 = {io_validin64_33,io_in64_33}; // @[Cat.scala 30:58]
  assign ingress2_8_io_in4_2 = {io_validin64_34,io_in64_34}; // @[Cat.scala 30:58]
  assign ingress2_8_io_in4_3 = {io_validin64_35,io_in64_35}; // @[Cat.scala 30:58]
  assign ingress2_8_io_ctrl = io_ctrl[63:56]; // @[BuildingBlock.scala 95:35]
  assign ingress2_9_clock = clock;
  assign ingress2_9_io_in4_0 = {io_validin64_36,io_in64_36}; // @[Cat.scala 30:58]
  assign ingress2_9_io_in4_1 = {io_validin64_37,io_in64_37}; // @[Cat.scala 30:58]
  assign ingress2_9_io_in4_2 = {io_validin64_38,io_in64_38}; // @[Cat.scala 30:58]
  assign ingress2_9_io_in4_3 = {io_validin64_39,io_in64_39}; // @[Cat.scala 30:58]
  assign ingress2_9_io_ctrl = io_ctrl[55:48]; // @[BuildingBlock.scala 95:35]
  assign ingress2_10_clock = clock;
  assign ingress2_10_io_in4_0 = {io_validin64_40,io_in64_40}; // @[Cat.scala 30:58]
  assign ingress2_10_io_in4_1 = {io_validin64_41,io_in64_41}; // @[Cat.scala 30:58]
  assign ingress2_10_io_in4_2 = {io_validin64_42,io_in64_42}; // @[Cat.scala 30:58]
  assign ingress2_10_io_in4_3 = {io_validin64_43,io_in64_43}; // @[Cat.scala 30:58]
  assign ingress2_10_io_ctrl = io_ctrl[47:40]; // @[BuildingBlock.scala 95:35]
  assign ingress2_11_clock = clock;
  assign ingress2_11_io_in4_0 = {io_validin64_44,io_in64_44}; // @[Cat.scala 30:58]
  assign ingress2_11_io_in4_1 = {io_validin64_45,io_in64_45}; // @[Cat.scala 30:58]
  assign ingress2_11_io_in4_2 = {io_validin64_46,io_in64_46}; // @[Cat.scala 30:58]
  assign ingress2_11_io_in4_3 = {io_validin64_47,io_in64_47}; // @[Cat.scala 30:58]
  assign ingress2_11_io_ctrl = io_ctrl[39:32]; // @[BuildingBlock.scala 95:35]
  assign ingress2_12_clock = clock;
  assign ingress2_12_io_in4_0 = {io_validin64_48,io_in64_48}; // @[Cat.scala 30:58]
  assign ingress2_12_io_in4_1 = {io_validin64_49,io_in64_49}; // @[Cat.scala 30:58]
  assign ingress2_12_io_in4_2 = {io_validin64_50,io_in64_50}; // @[Cat.scala 30:58]
  assign ingress2_12_io_in4_3 = {io_validin64_51,io_in64_51}; // @[Cat.scala 30:58]
  assign ingress2_12_io_ctrl = io_ctrl[31:24]; // @[BuildingBlock.scala 95:35]
  assign ingress2_13_clock = clock;
  assign ingress2_13_io_in4_0 = {io_validin64_52,io_in64_52}; // @[Cat.scala 30:58]
  assign ingress2_13_io_in4_1 = {io_validin64_53,io_in64_53}; // @[Cat.scala 30:58]
  assign ingress2_13_io_in4_2 = {io_validin64_54,io_in64_54}; // @[Cat.scala 30:58]
  assign ingress2_13_io_in4_3 = {io_validin64_55,io_in64_55}; // @[Cat.scala 30:58]
  assign ingress2_13_io_ctrl = io_ctrl[23:16]; // @[BuildingBlock.scala 95:35]
  assign ingress2_14_clock = clock;
  assign ingress2_14_io_in4_0 = {io_validin64_56,io_in64_56}; // @[Cat.scala 30:58]
  assign ingress2_14_io_in4_1 = {io_validin64_57,io_in64_57}; // @[Cat.scala 30:58]
  assign ingress2_14_io_in4_2 = {io_validin64_58,io_in64_58}; // @[Cat.scala 30:58]
  assign ingress2_14_io_in4_3 = {io_validin64_59,io_in64_59}; // @[Cat.scala 30:58]
  assign ingress2_14_io_ctrl = io_ctrl[15:8]; // @[BuildingBlock.scala 95:35]
  assign ingress2_15_clock = clock;
  assign ingress2_15_io_in4_0 = {io_validin64_60,io_in64_60}; // @[Cat.scala 30:58]
  assign ingress2_15_io_in4_1 = {io_validin64_61,io_in64_61}; // @[Cat.scala 30:58]
  assign ingress2_15_io_in4_2 = {io_validin64_62,io_in64_62}; // @[Cat.scala 30:58]
  assign ingress2_15_io_in4_3 = {io_validin64_63,io_in64_63}; // @[Cat.scala 30:58]
  assign ingress2_15_io_ctrl = io_ctrl[7:0]; // @[BuildingBlock.scala 95:35]
  always @(posedge clock) begin
    tag_Tag <= io_tagin_Tag; // @[BuildingBlock.scala 76:20]
    tag_RoundCnt <= io_tagin_RoundCnt; // @[BuildingBlock.scala 76:20]
    addr <= io_addrin; // @[BuildingBlock.scala 78:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_Tag = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  tag_RoundCnt = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  addr = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CLOSegress1(
  input          clock,
  input  [63:0]  io_in64_0,
  input  [63:0]  io_in64_1,
  input  [63:0]  io_in64_2,
  input  [63:0]  io_in64_3,
  input  [63:0]  io_in64_4,
  input  [63:0]  io_in64_5,
  input  [63:0]  io_in64_6,
  input  [63:0]  io_in64_7,
  input  [63:0]  io_in64_8,
  input  [63:0]  io_in64_9,
  input  [63:0]  io_in64_10,
  input  [63:0]  io_in64_11,
  input  [63:0]  io_in64_12,
  input  [63:0]  io_in64_13,
  input  [63:0]  io_in64_14,
  input  [63:0]  io_in64_15,
  input  [63:0]  io_in64_16,
  input  [63:0]  io_in64_17,
  input  [63:0]  io_in64_18,
  input  [63:0]  io_in64_19,
  input  [63:0]  io_in64_20,
  input  [63:0]  io_in64_21,
  input  [63:0]  io_in64_22,
  input  [63:0]  io_in64_23,
  input  [63:0]  io_in64_24,
  input  [63:0]  io_in64_25,
  input  [63:0]  io_in64_26,
  input  [63:0]  io_in64_27,
  input  [63:0]  io_in64_28,
  input  [63:0]  io_in64_29,
  input  [63:0]  io_in64_30,
  input  [63:0]  io_in64_31,
  input  [63:0]  io_in64_32,
  input  [63:0]  io_in64_33,
  input  [63:0]  io_in64_34,
  input  [63:0]  io_in64_35,
  input  [63:0]  io_in64_36,
  input  [63:0]  io_in64_37,
  input  [63:0]  io_in64_38,
  input  [63:0]  io_in64_39,
  input  [63:0]  io_in64_40,
  input  [63:0]  io_in64_41,
  input  [63:0]  io_in64_42,
  input  [63:0]  io_in64_43,
  input  [63:0]  io_in64_44,
  input  [63:0]  io_in64_45,
  input  [63:0]  io_in64_46,
  input  [63:0]  io_in64_47,
  input  [63:0]  io_in64_48,
  input  [63:0]  io_in64_49,
  input  [63:0]  io_in64_50,
  input  [63:0]  io_in64_51,
  input  [63:0]  io_in64_52,
  input  [63:0]  io_in64_53,
  input  [63:0]  io_in64_54,
  input  [63:0]  io_in64_55,
  input  [63:0]  io_in64_56,
  input  [63:0]  io_in64_57,
  input  [63:0]  io_in64_58,
  input  [63:0]  io_in64_59,
  input  [63:0]  io_in64_60,
  input  [63:0]  io_in64_61,
  input  [63:0]  io_in64_62,
  input  [63:0]  io_in64_63,
  input          io_validin64_0,
  input          io_validin64_1,
  input          io_validin64_2,
  input          io_validin64_3,
  input          io_validin64_4,
  input          io_validin64_5,
  input          io_validin64_6,
  input          io_validin64_7,
  input          io_validin64_8,
  input          io_validin64_9,
  input          io_validin64_10,
  input          io_validin64_11,
  input          io_validin64_12,
  input          io_validin64_13,
  input          io_validin64_14,
  input          io_validin64_15,
  input          io_validin64_16,
  input          io_validin64_17,
  input          io_validin64_18,
  input          io_validin64_19,
  input          io_validin64_20,
  input          io_validin64_21,
  input          io_validin64_22,
  input          io_validin64_23,
  input          io_validin64_24,
  input          io_validin64_25,
  input          io_validin64_26,
  input          io_validin64_27,
  input          io_validin64_28,
  input          io_validin64_29,
  input          io_validin64_30,
  input          io_validin64_31,
  input          io_validin64_32,
  input          io_validin64_33,
  input          io_validin64_34,
  input          io_validin64_35,
  input          io_validin64_36,
  input          io_validin64_37,
  input          io_validin64_38,
  input          io_validin64_39,
  input          io_validin64_40,
  input          io_validin64_41,
  input          io_validin64_42,
  input          io_validin64_43,
  input          io_validin64_44,
  input          io_validin64_45,
  input          io_validin64_46,
  input          io_validin64_47,
  input          io_validin64_48,
  input          io_validin64_49,
  input          io_validin64_50,
  input          io_validin64_51,
  input          io_validin64_52,
  input          io_validin64_53,
  input          io_validin64_54,
  input          io_validin64_55,
  input          io_validin64_56,
  input          io_validin64_57,
  input          io_validin64_58,
  input          io_validin64_59,
  input          io_validin64_60,
  input          io_validin64_61,
  input          io_validin64_62,
  input          io_validin64_63,
  input  [1:0]   io_tagin_Tag,
  input  [2:0]   io_tagin_RoundCnt,
  input  [7:0]   io_addrin,
  output [63:0]  io_out64_0,
  output [63:0]  io_out64_1,
  output [63:0]  io_out64_2,
  output [63:0]  io_out64_3,
  output [63:0]  io_out64_4,
  output [63:0]  io_out64_5,
  output [63:0]  io_out64_6,
  output [63:0]  io_out64_7,
  output [63:0]  io_out64_8,
  output [63:0]  io_out64_9,
  output [63:0]  io_out64_10,
  output [63:0]  io_out64_11,
  output [63:0]  io_out64_12,
  output [63:0]  io_out64_13,
  output [63:0]  io_out64_14,
  output [63:0]  io_out64_15,
  output [63:0]  io_out64_16,
  output [63:0]  io_out64_17,
  output [63:0]  io_out64_18,
  output [63:0]  io_out64_19,
  output [63:0]  io_out64_20,
  output [63:0]  io_out64_21,
  output [63:0]  io_out64_22,
  output [63:0]  io_out64_23,
  output [63:0]  io_out64_24,
  output [63:0]  io_out64_25,
  output [63:0]  io_out64_26,
  output [63:0]  io_out64_27,
  output [63:0]  io_out64_28,
  output [63:0]  io_out64_29,
  output [63:0]  io_out64_30,
  output [63:0]  io_out64_31,
  output [63:0]  io_out64_32,
  output [63:0]  io_out64_33,
  output [63:0]  io_out64_34,
  output [63:0]  io_out64_35,
  output [63:0]  io_out64_36,
  output [63:0]  io_out64_37,
  output [63:0]  io_out64_38,
  output [63:0]  io_out64_39,
  output [63:0]  io_out64_40,
  output [63:0]  io_out64_41,
  output [63:0]  io_out64_42,
  output [63:0]  io_out64_43,
  output [63:0]  io_out64_44,
  output [63:0]  io_out64_45,
  output [63:0]  io_out64_46,
  output [63:0]  io_out64_47,
  output [63:0]  io_out64_48,
  output [63:0]  io_out64_49,
  output [63:0]  io_out64_50,
  output [63:0]  io_out64_51,
  output [63:0]  io_out64_52,
  output [63:0]  io_out64_53,
  output [63:0]  io_out64_54,
  output [63:0]  io_out64_55,
  output [63:0]  io_out64_56,
  output [63:0]  io_out64_57,
  output [63:0]  io_out64_58,
  output [63:0]  io_out64_59,
  output [63:0]  io_out64_60,
  output [63:0]  io_out64_61,
  output [63:0]  io_out64_62,
  output [63:0]  io_out64_63,
  output         io_validout64_0,
  output         io_validout64_1,
  output         io_validout64_2,
  output         io_validout64_3,
  output         io_validout64_4,
  output         io_validout64_5,
  output         io_validout64_6,
  output         io_validout64_7,
  output         io_validout64_8,
  output         io_validout64_9,
  output         io_validout64_10,
  output         io_validout64_11,
  output         io_validout64_12,
  output         io_validout64_13,
  output         io_validout64_14,
  output         io_validout64_15,
  output         io_validout64_16,
  output         io_validout64_17,
  output         io_validout64_18,
  output         io_validout64_19,
  output         io_validout64_20,
  output         io_validout64_21,
  output         io_validout64_22,
  output         io_validout64_23,
  output         io_validout64_24,
  output         io_validout64_25,
  output         io_validout64_26,
  output         io_validout64_27,
  output         io_validout64_28,
  output         io_validout64_29,
  output         io_validout64_30,
  output         io_validout64_31,
  output         io_validout64_32,
  output         io_validout64_33,
  output         io_validout64_34,
  output         io_validout64_35,
  output         io_validout64_36,
  output         io_validout64_37,
  output         io_validout64_38,
  output         io_validout64_39,
  output         io_validout64_40,
  output         io_validout64_41,
  output         io_validout64_42,
  output         io_validout64_43,
  output         io_validout64_44,
  output         io_validout64_45,
  output         io_validout64_46,
  output         io_validout64_47,
  output         io_validout64_48,
  output         io_validout64_49,
  output         io_validout64_50,
  output         io_validout64_51,
  output         io_validout64_52,
  output         io_validout64_53,
  output         io_validout64_54,
  output         io_validout64_55,
  output         io_validout64_56,
  output         io_validout64_57,
  output         io_validout64_58,
  output         io_validout64_59,
  output         io_validout64_60,
  output         io_validout64_61,
  output         io_validout64_62,
  output         io_validout64_63,
  output [1:0]   io_tagout_Tag,
  output [2:0]   io_tagout_RoundCnt,
  output [7:0]   io_addrout,
  input  [127:0] io_ctrl
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  egress1_0_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_0_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_0_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_0_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_0_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_0_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_0_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_0_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_0_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_0_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_1_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_1_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_1_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_1_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_1_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_1_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_1_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_1_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_1_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_1_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_2_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_2_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_2_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_2_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_2_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_2_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_2_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_2_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_2_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_2_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_3_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_3_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_3_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_3_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_3_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_3_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_3_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_3_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_3_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_3_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_4_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_4_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_4_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_4_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_4_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_4_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_4_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_4_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_4_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_4_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_5_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_5_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_5_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_5_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_5_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_5_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_5_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_5_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_5_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_5_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_6_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_6_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_6_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_6_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_6_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_6_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_6_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_6_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_6_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_6_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_7_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_7_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_7_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_7_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_7_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_7_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_7_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_7_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_7_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_7_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_8_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_8_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_8_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_8_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_8_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_8_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_8_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_8_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_8_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_8_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_9_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_9_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_9_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_9_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_9_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_9_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_9_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_9_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_9_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_9_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_10_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_10_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_10_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_10_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_10_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_10_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_10_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_10_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_10_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_10_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_11_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_11_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_11_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_11_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_11_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_11_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_11_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_11_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_11_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_11_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_12_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_12_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_12_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_12_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_12_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_12_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_12_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_12_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_12_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_12_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_13_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_13_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_13_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_13_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_13_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_13_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_13_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_13_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_13_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_13_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_14_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_14_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_14_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_14_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_14_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_14_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_14_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_14_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_14_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_14_io_ctrl; // @[BuildingBlock.scala 148:51]
  wire  egress1_15_clock; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_15_io_in4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_15_io_in4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_15_io_in4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_15_io_in4_3; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_15_io_out4_0; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_15_io_out4_1; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_15_io_out4_2; // @[BuildingBlock.scala 148:51]
  wire [64:0] egress1_15_io_out4_3; // @[BuildingBlock.scala 148:51]
  wire [7:0] egress1_15_io_ctrl; // @[BuildingBlock.scala 148:51]
  reg [1:0] tag_Tag; // @[BuildingBlock.scala 149:20]
  reg [2:0] tag_RoundCnt; // @[BuildingBlock.scala 149:20]
  reg [7:0] addr; // @[BuildingBlock.scala 151:21]
  CLOScell4 egress1_0 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_0_clock),
    .io_in4_0(egress1_0_io_in4_0),
    .io_in4_1(egress1_0_io_in4_1),
    .io_in4_2(egress1_0_io_in4_2),
    .io_in4_3(egress1_0_io_in4_3),
    .io_out4_0(egress1_0_io_out4_0),
    .io_out4_1(egress1_0_io_out4_1),
    .io_out4_2(egress1_0_io_out4_2),
    .io_out4_3(egress1_0_io_out4_3),
    .io_ctrl(egress1_0_io_ctrl)
  );
  CLOScell4 egress1_1 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_1_clock),
    .io_in4_0(egress1_1_io_in4_0),
    .io_in4_1(egress1_1_io_in4_1),
    .io_in4_2(egress1_1_io_in4_2),
    .io_in4_3(egress1_1_io_in4_3),
    .io_out4_0(egress1_1_io_out4_0),
    .io_out4_1(egress1_1_io_out4_1),
    .io_out4_2(egress1_1_io_out4_2),
    .io_out4_3(egress1_1_io_out4_3),
    .io_ctrl(egress1_1_io_ctrl)
  );
  CLOScell4 egress1_2 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_2_clock),
    .io_in4_0(egress1_2_io_in4_0),
    .io_in4_1(egress1_2_io_in4_1),
    .io_in4_2(egress1_2_io_in4_2),
    .io_in4_3(egress1_2_io_in4_3),
    .io_out4_0(egress1_2_io_out4_0),
    .io_out4_1(egress1_2_io_out4_1),
    .io_out4_2(egress1_2_io_out4_2),
    .io_out4_3(egress1_2_io_out4_3),
    .io_ctrl(egress1_2_io_ctrl)
  );
  CLOScell4 egress1_3 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_3_clock),
    .io_in4_0(egress1_3_io_in4_0),
    .io_in4_1(egress1_3_io_in4_1),
    .io_in4_2(egress1_3_io_in4_2),
    .io_in4_3(egress1_3_io_in4_3),
    .io_out4_0(egress1_3_io_out4_0),
    .io_out4_1(egress1_3_io_out4_1),
    .io_out4_2(egress1_3_io_out4_2),
    .io_out4_3(egress1_3_io_out4_3),
    .io_ctrl(egress1_3_io_ctrl)
  );
  CLOScell4 egress1_4 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_4_clock),
    .io_in4_0(egress1_4_io_in4_0),
    .io_in4_1(egress1_4_io_in4_1),
    .io_in4_2(egress1_4_io_in4_2),
    .io_in4_3(egress1_4_io_in4_3),
    .io_out4_0(egress1_4_io_out4_0),
    .io_out4_1(egress1_4_io_out4_1),
    .io_out4_2(egress1_4_io_out4_2),
    .io_out4_3(egress1_4_io_out4_3),
    .io_ctrl(egress1_4_io_ctrl)
  );
  CLOScell4 egress1_5 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_5_clock),
    .io_in4_0(egress1_5_io_in4_0),
    .io_in4_1(egress1_5_io_in4_1),
    .io_in4_2(egress1_5_io_in4_2),
    .io_in4_3(egress1_5_io_in4_3),
    .io_out4_0(egress1_5_io_out4_0),
    .io_out4_1(egress1_5_io_out4_1),
    .io_out4_2(egress1_5_io_out4_2),
    .io_out4_3(egress1_5_io_out4_3),
    .io_ctrl(egress1_5_io_ctrl)
  );
  CLOScell4 egress1_6 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_6_clock),
    .io_in4_0(egress1_6_io_in4_0),
    .io_in4_1(egress1_6_io_in4_1),
    .io_in4_2(egress1_6_io_in4_2),
    .io_in4_3(egress1_6_io_in4_3),
    .io_out4_0(egress1_6_io_out4_0),
    .io_out4_1(egress1_6_io_out4_1),
    .io_out4_2(egress1_6_io_out4_2),
    .io_out4_3(egress1_6_io_out4_3),
    .io_ctrl(egress1_6_io_ctrl)
  );
  CLOScell4 egress1_7 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_7_clock),
    .io_in4_0(egress1_7_io_in4_0),
    .io_in4_1(egress1_7_io_in4_1),
    .io_in4_2(egress1_7_io_in4_2),
    .io_in4_3(egress1_7_io_in4_3),
    .io_out4_0(egress1_7_io_out4_0),
    .io_out4_1(egress1_7_io_out4_1),
    .io_out4_2(egress1_7_io_out4_2),
    .io_out4_3(egress1_7_io_out4_3),
    .io_ctrl(egress1_7_io_ctrl)
  );
  CLOScell4 egress1_8 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_8_clock),
    .io_in4_0(egress1_8_io_in4_0),
    .io_in4_1(egress1_8_io_in4_1),
    .io_in4_2(egress1_8_io_in4_2),
    .io_in4_3(egress1_8_io_in4_3),
    .io_out4_0(egress1_8_io_out4_0),
    .io_out4_1(egress1_8_io_out4_1),
    .io_out4_2(egress1_8_io_out4_2),
    .io_out4_3(egress1_8_io_out4_3),
    .io_ctrl(egress1_8_io_ctrl)
  );
  CLOScell4 egress1_9 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_9_clock),
    .io_in4_0(egress1_9_io_in4_0),
    .io_in4_1(egress1_9_io_in4_1),
    .io_in4_2(egress1_9_io_in4_2),
    .io_in4_3(egress1_9_io_in4_3),
    .io_out4_0(egress1_9_io_out4_0),
    .io_out4_1(egress1_9_io_out4_1),
    .io_out4_2(egress1_9_io_out4_2),
    .io_out4_3(egress1_9_io_out4_3),
    .io_ctrl(egress1_9_io_ctrl)
  );
  CLOScell4 egress1_10 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_10_clock),
    .io_in4_0(egress1_10_io_in4_0),
    .io_in4_1(egress1_10_io_in4_1),
    .io_in4_2(egress1_10_io_in4_2),
    .io_in4_3(egress1_10_io_in4_3),
    .io_out4_0(egress1_10_io_out4_0),
    .io_out4_1(egress1_10_io_out4_1),
    .io_out4_2(egress1_10_io_out4_2),
    .io_out4_3(egress1_10_io_out4_3),
    .io_ctrl(egress1_10_io_ctrl)
  );
  CLOScell4 egress1_11 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_11_clock),
    .io_in4_0(egress1_11_io_in4_0),
    .io_in4_1(egress1_11_io_in4_1),
    .io_in4_2(egress1_11_io_in4_2),
    .io_in4_3(egress1_11_io_in4_3),
    .io_out4_0(egress1_11_io_out4_0),
    .io_out4_1(egress1_11_io_out4_1),
    .io_out4_2(egress1_11_io_out4_2),
    .io_out4_3(egress1_11_io_out4_3),
    .io_ctrl(egress1_11_io_ctrl)
  );
  CLOScell4 egress1_12 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_12_clock),
    .io_in4_0(egress1_12_io_in4_0),
    .io_in4_1(egress1_12_io_in4_1),
    .io_in4_2(egress1_12_io_in4_2),
    .io_in4_3(egress1_12_io_in4_3),
    .io_out4_0(egress1_12_io_out4_0),
    .io_out4_1(egress1_12_io_out4_1),
    .io_out4_2(egress1_12_io_out4_2),
    .io_out4_3(egress1_12_io_out4_3),
    .io_ctrl(egress1_12_io_ctrl)
  );
  CLOScell4 egress1_13 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_13_clock),
    .io_in4_0(egress1_13_io_in4_0),
    .io_in4_1(egress1_13_io_in4_1),
    .io_in4_2(egress1_13_io_in4_2),
    .io_in4_3(egress1_13_io_in4_3),
    .io_out4_0(egress1_13_io_out4_0),
    .io_out4_1(egress1_13_io_out4_1),
    .io_out4_2(egress1_13_io_out4_2),
    .io_out4_3(egress1_13_io_out4_3),
    .io_ctrl(egress1_13_io_ctrl)
  );
  CLOScell4 egress1_14 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_14_clock),
    .io_in4_0(egress1_14_io_in4_0),
    .io_in4_1(egress1_14_io_in4_1),
    .io_in4_2(egress1_14_io_in4_2),
    .io_in4_3(egress1_14_io_in4_3),
    .io_out4_0(egress1_14_io_out4_0),
    .io_out4_1(egress1_14_io_out4_1),
    .io_out4_2(egress1_14_io_out4_2),
    .io_out4_3(egress1_14_io_out4_3),
    .io_ctrl(egress1_14_io_ctrl)
  );
  CLOScell4 egress1_15 ( // @[BuildingBlock.scala 148:51]
    .clock(egress1_15_clock),
    .io_in4_0(egress1_15_io_in4_0),
    .io_in4_1(egress1_15_io_in4_1),
    .io_in4_2(egress1_15_io_in4_2),
    .io_in4_3(egress1_15_io_in4_3),
    .io_out4_0(egress1_15_io_out4_0),
    .io_out4_1(egress1_15_io_out4_1),
    .io_out4_2(egress1_15_io_out4_2),
    .io_out4_3(egress1_15_io_out4_3),
    .io_ctrl(egress1_15_io_ctrl)
  );
  assign io_out64_0 = egress1_0_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_1 = egress1_4_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_2 = egress1_8_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_3 = egress1_12_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_4 = egress1_0_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_5 = egress1_4_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_6 = egress1_8_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_7 = egress1_12_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_8 = egress1_0_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_9 = egress1_4_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_10 = egress1_8_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_11 = egress1_12_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_12 = egress1_0_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_13 = egress1_4_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_14 = egress1_8_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_15 = egress1_12_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_16 = egress1_1_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_17 = egress1_5_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_18 = egress1_9_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_19 = egress1_13_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_20 = egress1_1_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_21 = egress1_5_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_22 = egress1_9_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_23 = egress1_13_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_24 = egress1_1_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_25 = egress1_5_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_26 = egress1_9_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_27 = egress1_13_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_28 = egress1_1_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_29 = egress1_5_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_30 = egress1_9_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_31 = egress1_13_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_32 = egress1_2_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_33 = egress1_6_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_34 = egress1_10_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_35 = egress1_14_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_36 = egress1_2_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_37 = egress1_6_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_38 = egress1_10_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_39 = egress1_14_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_40 = egress1_2_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_41 = egress1_6_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_42 = egress1_10_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_43 = egress1_14_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_44 = egress1_2_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_45 = egress1_6_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_46 = egress1_10_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_47 = egress1_14_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_48 = egress1_3_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_49 = egress1_7_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_50 = egress1_11_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_51 = egress1_15_io_out4_0[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_52 = egress1_3_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_53 = egress1_7_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_54 = egress1_11_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_55 = egress1_15_io_out4_1[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_56 = egress1_3_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_57 = egress1_7_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_58 = egress1_11_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_59 = egress1_15_io_out4_2[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_60 = egress1_3_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_61 = egress1_7_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_62 = egress1_11_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_out64_63 = egress1_15_io_out4_3[63:0]; // @[BuildingBlock.scala 170:58]
  assign io_validout64_0 = egress1_0_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_1 = egress1_4_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_2 = egress1_8_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_3 = egress1_12_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_4 = egress1_0_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_5 = egress1_4_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_6 = egress1_8_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_7 = egress1_12_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_8 = egress1_0_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_9 = egress1_4_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_10 = egress1_8_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_11 = egress1_12_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_12 = egress1_0_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_13 = egress1_4_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_14 = egress1_8_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_15 = egress1_12_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_16 = egress1_1_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_17 = egress1_5_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_18 = egress1_9_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_19 = egress1_13_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_20 = egress1_1_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_21 = egress1_5_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_22 = egress1_9_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_23 = egress1_13_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_24 = egress1_1_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_25 = egress1_5_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_26 = egress1_9_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_27 = egress1_13_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_28 = egress1_1_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_29 = egress1_5_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_30 = egress1_9_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_31 = egress1_13_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_32 = egress1_2_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_33 = egress1_6_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_34 = egress1_10_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_35 = egress1_14_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_36 = egress1_2_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_37 = egress1_6_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_38 = egress1_10_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_39 = egress1_14_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_40 = egress1_2_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_41 = egress1_6_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_42 = egress1_10_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_43 = egress1_14_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_44 = egress1_2_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_45 = egress1_6_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_46 = egress1_10_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_47 = egress1_14_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_48 = egress1_3_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_49 = egress1_7_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_50 = egress1_11_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_51 = egress1_15_io_out4_0[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_52 = egress1_3_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_53 = egress1_7_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_54 = egress1_11_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_55 = egress1_15_io_out4_1[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_56 = egress1_3_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_57 = egress1_7_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_58 = egress1_11_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_59 = egress1_15_io_out4_2[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_60 = egress1_3_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_61 = egress1_7_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_62 = egress1_11_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_validout64_63 = egress1_15_io_out4_3[64]; // @[BuildingBlock.scala 171:63]
  assign io_tagout_Tag = tag_Tag; // @[BuildingBlock.scala 150:13]
  assign io_tagout_RoundCnt = tag_RoundCnt; // @[BuildingBlock.scala 150:13]
  assign io_addrout = addr; // @[BuildingBlock.scala 152:14]
  assign egress1_0_clock = clock;
  assign egress1_0_io_in4_0 = {io_validin64_0,io_in64_0}; // @[Cat.scala 30:58]
  assign egress1_0_io_in4_1 = {io_validin64_1,io_in64_1}; // @[Cat.scala 30:58]
  assign egress1_0_io_in4_2 = {io_validin64_2,io_in64_2}; // @[Cat.scala 30:58]
  assign egress1_0_io_in4_3 = {io_validin64_3,io_in64_3}; // @[Cat.scala 30:58]
  assign egress1_0_io_ctrl = io_ctrl[127:120]; // @[BuildingBlock.scala 177:34]
  assign egress1_1_clock = clock;
  assign egress1_1_io_in4_0 = {io_validin64_4,io_in64_4}; // @[Cat.scala 30:58]
  assign egress1_1_io_in4_1 = {io_validin64_5,io_in64_5}; // @[Cat.scala 30:58]
  assign egress1_1_io_in4_2 = {io_validin64_6,io_in64_6}; // @[Cat.scala 30:58]
  assign egress1_1_io_in4_3 = {io_validin64_7,io_in64_7}; // @[Cat.scala 30:58]
  assign egress1_1_io_ctrl = io_ctrl[119:112]; // @[BuildingBlock.scala 177:34]
  assign egress1_2_clock = clock;
  assign egress1_2_io_in4_0 = {io_validin64_8,io_in64_8}; // @[Cat.scala 30:58]
  assign egress1_2_io_in4_1 = {io_validin64_9,io_in64_9}; // @[Cat.scala 30:58]
  assign egress1_2_io_in4_2 = {io_validin64_10,io_in64_10}; // @[Cat.scala 30:58]
  assign egress1_2_io_in4_3 = {io_validin64_11,io_in64_11}; // @[Cat.scala 30:58]
  assign egress1_2_io_ctrl = io_ctrl[111:104]; // @[BuildingBlock.scala 177:34]
  assign egress1_3_clock = clock;
  assign egress1_3_io_in4_0 = {io_validin64_12,io_in64_12}; // @[Cat.scala 30:58]
  assign egress1_3_io_in4_1 = {io_validin64_13,io_in64_13}; // @[Cat.scala 30:58]
  assign egress1_3_io_in4_2 = {io_validin64_14,io_in64_14}; // @[Cat.scala 30:58]
  assign egress1_3_io_in4_3 = {io_validin64_15,io_in64_15}; // @[Cat.scala 30:58]
  assign egress1_3_io_ctrl = io_ctrl[103:96]; // @[BuildingBlock.scala 177:34]
  assign egress1_4_clock = clock;
  assign egress1_4_io_in4_0 = {io_validin64_16,io_in64_16}; // @[Cat.scala 30:58]
  assign egress1_4_io_in4_1 = {io_validin64_17,io_in64_17}; // @[Cat.scala 30:58]
  assign egress1_4_io_in4_2 = {io_validin64_18,io_in64_18}; // @[Cat.scala 30:58]
  assign egress1_4_io_in4_3 = {io_validin64_19,io_in64_19}; // @[Cat.scala 30:58]
  assign egress1_4_io_ctrl = io_ctrl[95:88]; // @[BuildingBlock.scala 177:34]
  assign egress1_5_clock = clock;
  assign egress1_5_io_in4_0 = {io_validin64_20,io_in64_20}; // @[Cat.scala 30:58]
  assign egress1_5_io_in4_1 = {io_validin64_21,io_in64_21}; // @[Cat.scala 30:58]
  assign egress1_5_io_in4_2 = {io_validin64_22,io_in64_22}; // @[Cat.scala 30:58]
  assign egress1_5_io_in4_3 = {io_validin64_23,io_in64_23}; // @[Cat.scala 30:58]
  assign egress1_5_io_ctrl = io_ctrl[87:80]; // @[BuildingBlock.scala 177:34]
  assign egress1_6_clock = clock;
  assign egress1_6_io_in4_0 = {io_validin64_24,io_in64_24}; // @[Cat.scala 30:58]
  assign egress1_6_io_in4_1 = {io_validin64_25,io_in64_25}; // @[Cat.scala 30:58]
  assign egress1_6_io_in4_2 = {io_validin64_26,io_in64_26}; // @[Cat.scala 30:58]
  assign egress1_6_io_in4_3 = {io_validin64_27,io_in64_27}; // @[Cat.scala 30:58]
  assign egress1_6_io_ctrl = io_ctrl[79:72]; // @[BuildingBlock.scala 177:34]
  assign egress1_7_clock = clock;
  assign egress1_7_io_in4_0 = {io_validin64_28,io_in64_28}; // @[Cat.scala 30:58]
  assign egress1_7_io_in4_1 = {io_validin64_29,io_in64_29}; // @[Cat.scala 30:58]
  assign egress1_7_io_in4_2 = {io_validin64_30,io_in64_30}; // @[Cat.scala 30:58]
  assign egress1_7_io_in4_3 = {io_validin64_31,io_in64_31}; // @[Cat.scala 30:58]
  assign egress1_7_io_ctrl = io_ctrl[71:64]; // @[BuildingBlock.scala 177:34]
  assign egress1_8_clock = clock;
  assign egress1_8_io_in4_0 = {io_validin64_32,io_in64_32}; // @[Cat.scala 30:58]
  assign egress1_8_io_in4_1 = {io_validin64_33,io_in64_33}; // @[Cat.scala 30:58]
  assign egress1_8_io_in4_2 = {io_validin64_34,io_in64_34}; // @[Cat.scala 30:58]
  assign egress1_8_io_in4_3 = {io_validin64_35,io_in64_35}; // @[Cat.scala 30:58]
  assign egress1_8_io_ctrl = io_ctrl[63:56]; // @[BuildingBlock.scala 177:34]
  assign egress1_9_clock = clock;
  assign egress1_9_io_in4_0 = {io_validin64_36,io_in64_36}; // @[Cat.scala 30:58]
  assign egress1_9_io_in4_1 = {io_validin64_37,io_in64_37}; // @[Cat.scala 30:58]
  assign egress1_9_io_in4_2 = {io_validin64_38,io_in64_38}; // @[Cat.scala 30:58]
  assign egress1_9_io_in4_3 = {io_validin64_39,io_in64_39}; // @[Cat.scala 30:58]
  assign egress1_9_io_ctrl = io_ctrl[55:48]; // @[BuildingBlock.scala 177:34]
  assign egress1_10_clock = clock;
  assign egress1_10_io_in4_0 = {io_validin64_40,io_in64_40}; // @[Cat.scala 30:58]
  assign egress1_10_io_in4_1 = {io_validin64_41,io_in64_41}; // @[Cat.scala 30:58]
  assign egress1_10_io_in4_2 = {io_validin64_42,io_in64_42}; // @[Cat.scala 30:58]
  assign egress1_10_io_in4_3 = {io_validin64_43,io_in64_43}; // @[Cat.scala 30:58]
  assign egress1_10_io_ctrl = io_ctrl[47:40]; // @[BuildingBlock.scala 177:34]
  assign egress1_11_clock = clock;
  assign egress1_11_io_in4_0 = {io_validin64_44,io_in64_44}; // @[Cat.scala 30:58]
  assign egress1_11_io_in4_1 = {io_validin64_45,io_in64_45}; // @[Cat.scala 30:58]
  assign egress1_11_io_in4_2 = {io_validin64_46,io_in64_46}; // @[Cat.scala 30:58]
  assign egress1_11_io_in4_3 = {io_validin64_47,io_in64_47}; // @[Cat.scala 30:58]
  assign egress1_11_io_ctrl = io_ctrl[39:32]; // @[BuildingBlock.scala 177:34]
  assign egress1_12_clock = clock;
  assign egress1_12_io_in4_0 = {io_validin64_48,io_in64_48}; // @[Cat.scala 30:58]
  assign egress1_12_io_in4_1 = {io_validin64_49,io_in64_49}; // @[Cat.scala 30:58]
  assign egress1_12_io_in4_2 = {io_validin64_50,io_in64_50}; // @[Cat.scala 30:58]
  assign egress1_12_io_in4_3 = {io_validin64_51,io_in64_51}; // @[Cat.scala 30:58]
  assign egress1_12_io_ctrl = io_ctrl[31:24]; // @[BuildingBlock.scala 177:34]
  assign egress1_13_clock = clock;
  assign egress1_13_io_in4_0 = {io_validin64_52,io_in64_52}; // @[Cat.scala 30:58]
  assign egress1_13_io_in4_1 = {io_validin64_53,io_in64_53}; // @[Cat.scala 30:58]
  assign egress1_13_io_in4_2 = {io_validin64_54,io_in64_54}; // @[Cat.scala 30:58]
  assign egress1_13_io_in4_3 = {io_validin64_55,io_in64_55}; // @[Cat.scala 30:58]
  assign egress1_13_io_ctrl = io_ctrl[23:16]; // @[BuildingBlock.scala 177:34]
  assign egress1_14_clock = clock;
  assign egress1_14_io_in4_0 = {io_validin64_56,io_in64_56}; // @[Cat.scala 30:58]
  assign egress1_14_io_in4_1 = {io_validin64_57,io_in64_57}; // @[Cat.scala 30:58]
  assign egress1_14_io_in4_2 = {io_validin64_58,io_in64_58}; // @[Cat.scala 30:58]
  assign egress1_14_io_in4_3 = {io_validin64_59,io_in64_59}; // @[Cat.scala 30:58]
  assign egress1_14_io_ctrl = io_ctrl[15:8]; // @[BuildingBlock.scala 177:34]
  assign egress1_15_clock = clock;
  assign egress1_15_io_in4_0 = {io_validin64_60,io_in64_60}; // @[Cat.scala 30:58]
  assign egress1_15_io_in4_1 = {io_validin64_61,io_in64_61}; // @[Cat.scala 30:58]
  assign egress1_15_io_in4_2 = {io_validin64_62,io_in64_62}; // @[Cat.scala 30:58]
  assign egress1_15_io_in4_3 = {io_validin64_63,io_in64_63}; // @[Cat.scala 30:58]
  assign egress1_15_io_ctrl = io_ctrl[7:0]; // @[BuildingBlock.scala 177:34]
  always @(posedge clock) begin
    tag_Tag <= io_tagin_Tag; // @[BuildingBlock.scala 149:20]
    tag_RoundCnt <= io_tagin_RoundCnt; // @[BuildingBlock.scala 149:20]
    addr <= io_addrin; // @[BuildingBlock.scala 151:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_Tag = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  tag_RoundCnt = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  addr = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CLOSegress2(
  input          clock,
  input  [63:0]  io_in64_0,
  input  [63:0]  io_in64_1,
  input  [63:0]  io_in64_2,
  input  [63:0]  io_in64_3,
  input  [63:0]  io_in64_4,
  input  [63:0]  io_in64_5,
  input  [63:0]  io_in64_6,
  input  [63:0]  io_in64_7,
  input  [63:0]  io_in64_8,
  input  [63:0]  io_in64_9,
  input  [63:0]  io_in64_10,
  input  [63:0]  io_in64_11,
  input  [63:0]  io_in64_12,
  input  [63:0]  io_in64_13,
  input  [63:0]  io_in64_14,
  input  [63:0]  io_in64_15,
  input  [63:0]  io_in64_16,
  input  [63:0]  io_in64_17,
  input  [63:0]  io_in64_18,
  input  [63:0]  io_in64_19,
  input  [63:0]  io_in64_20,
  input  [63:0]  io_in64_21,
  input  [63:0]  io_in64_22,
  input  [63:0]  io_in64_23,
  input  [63:0]  io_in64_24,
  input  [63:0]  io_in64_25,
  input  [63:0]  io_in64_26,
  input  [63:0]  io_in64_27,
  input  [63:0]  io_in64_28,
  input  [63:0]  io_in64_29,
  input  [63:0]  io_in64_30,
  input  [63:0]  io_in64_31,
  input  [63:0]  io_in64_32,
  input  [63:0]  io_in64_33,
  input  [63:0]  io_in64_34,
  input  [63:0]  io_in64_35,
  input  [63:0]  io_in64_36,
  input  [63:0]  io_in64_37,
  input  [63:0]  io_in64_38,
  input  [63:0]  io_in64_39,
  input  [63:0]  io_in64_40,
  input  [63:0]  io_in64_41,
  input  [63:0]  io_in64_42,
  input  [63:0]  io_in64_43,
  input  [63:0]  io_in64_44,
  input  [63:0]  io_in64_45,
  input  [63:0]  io_in64_46,
  input  [63:0]  io_in64_47,
  input  [63:0]  io_in64_48,
  input  [63:0]  io_in64_49,
  input  [63:0]  io_in64_50,
  input  [63:0]  io_in64_51,
  input  [63:0]  io_in64_52,
  input  [63:0]  io_in64_53,
  input  [63:0]  io_in64_54,
  input  [63:0]  io_in64_55,
  input  [63:0]  io_in64_56,
  input  [63:0]  io_in64_57,
  input  [63:0]  io_in64_58,
  input  [63:0]  io_in64_59,
  input  [63:0]  io_in64_60,
  input  [63:0]  io_in64_61,
  input  [63:0]  io_in64_62,
  input  [63:0]  io_in64_63,
  input          io_validin64_0,
  input          io_validin64_1,
  input          io_validin64_2,
  input          io_validin64_3,
  input          io_validin64_4,
  input          io_validin64_5,
  input          io_validin64_6,
  input          io_validin64_7,
  input          io_validin64_8,
  input          io_validin64_9,
  input          io_validin64_10,
  input          io_validin64_11,
  input          io_validin64_12,
  input          io_validin64_13,
  input          io_validin64_14,
  input          io_validin64_15,
  input          io_validin64_16,
  input          io_validin64_17,
  input          io_validin64_18,
  input          io_validin64_19,
  input          io_validin64_20,
  input          io_validin64_21,
  input          io_validin64_22,
  input          io_validin64_23,
  input          io_validin64_24,
  input          io_validin64_25,
  input          io_validin64_26,
  input          io_validin64_27,
  input          io_validin64_28,
  input          io_validin64_29,
  input          io_validin64_30,
  input          io_validin64_31,
  input          io_validin64_32,
  input          io_validin64_33,
  input          io_validin64_34,
  input          io_validin64_35,
  input          io_validin64_36,
  input          io_validin64_37,
  input          io_validin64_38,
  input          io_validin64_39,
  input          io_validin64_40,
  input          io_validin64_41,
  input          io_validin64_42,
  input          io_validin64_43,
  input          io_validin64_44,
  input          io_validin64_45,
  input          io_validin64_46,
  input          io_validin64_47,
  input          io_validin64_48,
  input          io_validin64_49,
  input          io_validin64_50,
  input          io_validin64_51,
  input          io_validin64_52,
  input          io_validin64_53,
  input          io_validin64_54,
  input          io_validin64_55,
  input          io_validin64_56,
  input          io_validin64_57,
  input          io_validin64_58,
  input          io_validin64_59,
  input          io_validin64_60,
  input          io_validin64_61,
  input          io_validin64_62,
  input          io_validin64_63,
  input  [1:0]   io_tagin_Tag,
  input  [2:0]   io_tagin_RoundCnt,
  input  [7:0]   io_addrin,
  output [63:0]  io_out64_0,
  output [63:0]  io_out64_1,
  output [63:0]  io_out64_2,
  output [63:0]  io_out64_3,
  output [63:0]  io_out64_4,
  output [63:0]  io_out64_5,
  output [63:0]  io_out64_6,
  output [63:0]  io_out64_7,
  output [63:0]  io_out64_8,
  output [63:0]  io_out64_9,
  output [63:0]  io_out64_10,
  output [63:0]  io_out64_11,
  output [63:0]  io_out64_12,
  output [63:0]  io_out64_13,
  output [63:0]  io_out64_14,
  output [63:0]  io_out64_15,
  output [63:0]  io_out64_16,
  output [63:0]  io_out64_17,
  output [63:0]  io_out64_18,
  output [63:0]  io_out64_19,
  output [63:0]  io_out64_20,
  output [63:0]  io_out64_21,
  output [63:0]  io_out64_22,
  output [63:0]  io_out64_23,
  output [63:0]  io_out64_24,
  output [63:0]  io_out64_25,
  output [63:0]  io_out64_26,
  output [63:0]  io_out64_27,
  output [63:0]  io_out64_28,
  output [63:0]  io_out64_29,
  output [63:0]  io_out64_30,
  output [63:0]  io_out64_31,
  output [63:0]  io_out64_32,
  output [63:0]  io_out64_33,
  output [63:0]  io_out64_34,
  output [63:0]  io_out64_35,
  output [63:0]  io_out64_36,
  output [63:0]  io_out64_37,
  output [63:0]  io_out64_38,
  output [63:0]  io_out64_39,
  output [63:0]  io_out64_40,
  output [63:0]  io_out64_41,
  output [63:0]  io_out64_42,
  output [63:0]  io_out64_43,
  output [63:0]  io_out64_44,
  output [63:0]  io_out64_45,
  output [63:0]  io_out64_46,
  output [63:0]  io_out64_47,
  output [63:0]  io_out64_48,
  output [63:0]  io_out64_49,
  output [63:0]  io_out64_50,
  output [63:0]  io_out64_51,
  output [63:0]  io_out64_52,
  output [63:0]  io_out64_53,
  output [63:0]  io_out64_54,
  output [63:0]  io_out64_55,
  output [63:0]  io_out64_56,
  output [63:0]  io_out64_57,
  output [63:0]  io_out64_58,
  output [63:0]  io_out64_59,
  output [63:0]  io_out64_60,
  output [63:0]  io_out64_61,
  output [63:0]  io_out64_62,
  output [63:0]  io_out64_63,
  output         io_validout64_0,
  output         io_validout64_1,
  output         io_validout64_2,
  output         io_validout64_3,
  output         io_validout64_4,
  output         io_validout64_5,
  output         io_validout64_6,
  output         io_validout64_7,
  output         io_validout64_8,
  output         io_validout64_9,
  output         io_validout64_10,
  output         io_validout64_11,
  output         io_validout64_12,
  output         io_validout64_13,
  output         io_validout64_14,
  output         io_validout64_15,
  output         io_validout64_16,
  output         io_validout64_17,
  output         io_validout64_18,
  output         io_validout64_19,
  output         io_validout64_20,
  output         io_validout64_21,
  output         io_validout64_22,
  output         io_validout64_23,
  output         io_validout64_24,
  output         io_validout64_25,
  output         io_validout64_26,
  output         io_validout64_27,
  output         io_validout64_28,
  output         io_validout64_29,
  output         io_validout64_30,
  output         io_validout64_31,
  output         io_validout64_32,
  output         io_validout64_33,
  output         io_validout64_34,
  output         io_validout64_35,
  output         io_validout64_36,
  output         io_validout64_37,
  output         io_validout64_38,
  output         io_validout64_39,
  output         io_validout64_40,
  output         io_validout64_41,
  output         io_validout64_42,
  output         io_validout64_43,
  output         io_validout64_44,
  output         io_validout64_45,
  output         io_validout64_46,
  output         io_validout64_47,
  output         io_validout64_48,
  output         io_validout64_49,
  output         io_validout64_50,
  output         io_validout64_51,
  output         io_validout64_52,
  output         io_validout64_53,
  output         io_validout64_54,
  output         io_validout64_55,
  output         io_validout64_56,
  output         io_validout64_57,
  output         io_validout64_58,
  output         io_validout64_59,
  output         io_validout64_60,
  output         io_validout64_61,
  output         io_validout64_62,
  output         io_validout64_63,
  output [1:0]   io_tagout_Tag,
  output [2:0]   io_tagout_RoundCnt,
  output [7:0]   io_addrout,
  input  [127:0] io_ctrl
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  egress2_0_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_0_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_0_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_0_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_0_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_0_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_0_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_0_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_0_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_0_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_1_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_1_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_1_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_1_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_1_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_1_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_1_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_1_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_1_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_1_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_2_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_2_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_2_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_2_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_2_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_2_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_2_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_2_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_2_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_2_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_3_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_3_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_3_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_3_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_3_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_3_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_3_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_3_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_3_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_3_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_4_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_4_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_4_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_4_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_4_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_4_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_4_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_4_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_4_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_4_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_5_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_5_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_5_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_5_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_5_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_5_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_5_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_5_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_5_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_5_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_6_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_6_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_6_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_6_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_6_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_6_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_6_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_6_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_6_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_6_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_7_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_7_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_7_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_7_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_7_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_7_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_7_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_7_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_7_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_7_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_8_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_8_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_8_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_8_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_8_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_8_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_8_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_8_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_8_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_8_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_9_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_9_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_9_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_9_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_9_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_9_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_9_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_9_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_9_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_9_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_10_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_10_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_10_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_10_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_10_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_10_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_10_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_10_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_10_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_10_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_11_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_11_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_11_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_11_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_11_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_11_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_11_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_11_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_11_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_11_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_12_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_12_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_12_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_12_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_12_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_12_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_12_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_12_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_12_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_12_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_13_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_13_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_13_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_13_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_13_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_13_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_13_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_13_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_13_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_13_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_14_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_14_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_14_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_14_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_14_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_14_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_14_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_14_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_14_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_14_io_ctrl; // @[BuildingBlock.scala 193:51]
  wire  egress2_15_clock; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_15_io_in4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_15_io_in4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_15_io_in4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_15_io_in4_3; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_15_io_out4_0; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_15_io_out4_1; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_15_io_out4_2; // @[BuildingBlock.scala 193:51]
  wire [64:0] egress2_15_io_out4_3; // @[BuildingBlock.scala 193:51]
  wire [7:0] egress2_15_io_ctrl; // @[BuildingBlock.scala 193:51]
  reg [1:0] tag_Tag; // @[BuildingBlock.scala 194:20]
  reg [2:0] tag_RoundCnt; // @[BuildingBlock.scala 194:20]
  reg [7:0] addr; // @[BuildingBlock.scala 196:21]
  CLOScell4 egress2_0 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_0_clock),
    .io_in4_0(egress2_0_io_in4_0),
    .io_in4_1(egress2_0_io_in4_1),
    .io_in4_2(egress2_0_io_in4_2),
    .io_in4_3(egress2_0_io_in4_3),
    .io_out4_0(egress2_0_io_out4_0),
    .io_out4_1(egress2_0_io_out4_1),
    .io_out4_2(egress2_0_io_out4_2),
    .io_out4_3(egress2_0_io_out4_3),
    .io_ctrl(egress2_0_io_ctrl)
  );
  CLOScell4 egress2_1 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_1_clock),
    .io_in4_0(egress2_1_io_in4_0),
    .io_in4_1(egress2_1_io_in4_1),
    .io_in4_2(egress2_1_io_in4_2),
    .io_in4_3(egress2_1_io_in4_3),
    .io_out4_0(egress2_1_io_out4_0),
    .io_out4_1(egress2_1_io_out4_1),
    .io_out4_2(egress2_1_io_out4_2),
    .io_out4_3(egress2_1_io_out4_3),
    .io_ctrl(egress2_1_io_ctrl)
  );
  CLOScell4 egress2_2 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_2_clock),
    .io_in4_0(egress2_2_io_in4_0),
    .io_in4_1(egress2_2_io_in4_1),
    .io_in4_2(egress2_2_io_in4_2),
    .io_in4_3(egress2_2_io_in4_3),
    .io_out4_0(egress2_2_io_out4_0),
    .io_out4_1(egress2_2_io_out4_1),
    .io_out4_2(egress2_2_io_out4_2),
    .io_out4_3(egress2_2_io_out4_3),
    .io_ctrl(egress2_2_io_ctrl)
  );
  CLOScell4 egress2_3 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_3_clock),
    .io_in4_0(egress2_3_io_in4_0),
    .io_in4_1(egress2_3_io_in4_1),
    .io_in4_2(egress2_3_io_in4_2),
    .io_in4_3(egress2_3_io_in4_3),
    .io_out4_0(egress2_3_io_out4_0),
    .io_out4_1(egress2_3_io_out4_1),
    .io_out4_2(egress2_3_io_out4_2),
    .io_out4_3(egress2_3_io_out4_3),
    .io_ctrl(egress2_3_io_ctrl)
  );
  CLOScell4 egress2_4 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_4_clock),
    .io_in4_0(egress2_4_io_in4_0),
    .io_in4_1(egress2_4_io_in4_1),
    .io_in4_2(egress2_4_io_in4_2),
    .io_in4_3(egress2_4_io_in4_3),
    .io_out4_0(egress2_4_io_out4_0),
    .io_out4_1(egress2_4_io_out4_1),
    .io_out4_2(egress2_4_io_out4_2),
    .io_out4_3(egress2_4_io_out4_3),
    .io_ctrl(egress2_4_io_ctrl)
  );
  CLOScell4 egress2_5 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_5_clock),
    .io_in4_0(egress2_5_io_in4_0),
    .io_in4_1(egress2_5_io_in4_1),
    .io_in4_2(egress2_5_io_in4_2),
    .io_in4_3(egress2_5_io_in4_3),
    .io_out4_0(egress2_5_io_out4_0),
    .io_out4_1(egress2_5_io_out4_1),
    .io_out4_2(egress2_5_io_out4_2),
    .io_out4_3(egress2_5_io_out4_3),
    .io_ctrl(egress2_5_io_ctrl)
  );
  CLOScell4 egress2_6 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_6_clock),
    .io_in4_0(egress2_6_io_in4_0),
    .io_in4_1(egress2_6_io_in4_1),
    .io_in4_2(egress2_6_io_in4_2),
    .io_in4_3(egress2_6_io_in4_3),
    .io_out4_0(egress2_6_io_out4_0),
    .io_out4_1(egress2_6_io_out4_1),
    .io_out4_2(egress2_6_io_out4_2),
    .io_out4_3(egress2_6_io_out4_3),
    .io_ctrl(egress2_6_io_ctrl)
  );
  CLOScell4 egress2_7 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_7_clock),
    .io_in4_0(egress2_7_io_in4_0),
    .io_in4_1(egress2_7_io_in4_1),
    .io_in4_2(egress2_7_io_in4_2),
    .io_in4_3(egress2_7_io_in4_3),
    .io_out4_0(egress2_7_io_out4_0),
    .io_out4_1(egress2_7_io_out4_1),
    .io_out4_2(egress2_7_io_out4_2),
    .io_out4_3(egress2_7_io_out4_3),
    .io_ctrl(egress2_7_io_ctrl)
  );
  CLOScell4 egress2_8 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_8_clock),
    .io_in4_0(egress2_8_io_in4_0),
    .io_in4_1(egress2_8_io_in4_1),
    .io_in4_2(egress2_8_io_in4_2),
    .io_in4_3(egress2_8_io_in4_3),
    .io_out4_0(egress2_8_io_out4_0),
    .io_out4_1(egress2_8_io_out4_1),
    .io_out4_2(egress2_8_io_out4_2),
    .io_out4_3(egress2_8_io_out4_3),
    .io_ctrl(egress2_8_io_ctrl)
  );
  CLOScell4 egress2_9 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_9_clock),
    .io_in4_0(egress2_9_io_in4_0),
    .io_in4_1(egress2_9_io_in4_1),
    .io_in4_2(egress2_9_io_in4_2),
    .io_in4_3(egress2_9_io_in4_3),
    .io_out4_0(egress2_9_io_out4_0),
    .io_out4_1(egress2_9_io_out4_1),
    .io_out4_2(egress2_9_io_out4_2),
    .io_out4_3(egress2_9_io_out4_3),
    .io_ctrl(egress2_9_io_ctrl)
  );
  CLOScell4 egress2_10 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_10_clock),
    .io_in4_0(egress2_10_io_in4_0),
    .io_in4_1(egress2_10_io_in4_1),
    .io_in4_2(egress2_10_io_in4_2),
    .io_in4_3(egress2_10_io_in4_3),
    .io_out4_0(egress2_10_io_out4_0),
    .io_out4_1(egress2_10_io_out4_1),
    .io_out4_2(egress2_10_io_out4_2),
    .io_out4_3(egress2_10_io_out4_3),
    .io_ctrl(egress2_10_io_ctrl)
  );
  CLOScell4 egress2_11 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_11_clock),
    .io_in4_0(egress2_11_io_in4_0),
    .io_in4_1(egress2_11_io_in4_1),
    .io_in4_2(egress2_11_io_in4_2),
    .io_in4_3(egress2_11_io_in4_3),
    .io_out4_0(egress2_11_io_out4_0),
    .io_out4_1(egress2_11_io_out4_1),
    .io_out4_2(egress2_11_io_out4_2),
    .io_out4_3(egress2_11_io_out4_3),
    .io_ctrl(egress2_11_io_ctrl)
  );
  CLOScell4 egress2_12 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_12_clock),
    .io_in4_0(egress2_12_io_in4_0),
    .io_in4_1(egress2_12_io_in4_1),
    .io_in4_2(egress2_12_io_in4_2),
    .io_in4_3(egress2_12_io_in4_3),
    .io_out4_0(egress2_12_io_out4_0),
    .io_out4_1(egress2_12_io_out4_1),
    .io_out4_2(egress2_12_io_out4_2),
    .io_out4_3(egress2_12_io_out4_3),
    .io_ctrl(egress2_12_io_ctrl)
  );
  CLOScell4 egress2_13 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_13_clock),
    .io_in4_0(egress2_13_io_in4_0),
    .io_in4_1(egress2_13_io_in4_1),
    .io_in4_2(egress2_13_io_in4_2),
    .io_in4_3(egress2_13_io_in4_3),
    .io_out4_0(egress2_13_io_out4_0),
    .io_out4_1(egress2_13_io_out4_1),
    .io_out4_2(egress2_13_io_out4_2),
    .io_out4_3(egress2_13_io_out4_3),
    .io_ctrl(egress2_13_io_ctrl)
  );
  CLOScell4 egress2_14 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_14_clock),
    .io_in4_0(egress2_14_io_in4_0),
    .io_in4_1(egress2_14_io_in4_1),
    .io_in4_2(egress2_14_io_in4_2),
    .io_in4_3(egress2_14_io_in4_3),
    .io_out4_0(egress2_14_io_out4_0),
    .io_out4_1(egress2_14_io_out4_1),
    .io_out4_2(egress2_14_io_out4_2),
    .io_out4_3(egress2_14_io_out4_3),
    .io_ctrl(egress2_14_io_ctrl)
  );
  CLOScell4 egress2_15 ( // @[BuildingBlock.scala 193:51]
    .clock(egress2_15_clock),
    .io_in4_0(egress2_15_io_in4_0),
    .io_in4_1(egress2_15_io_in4_1),
    .io_in4_2(egress2_15_io_in4_2),
    .io_in4_3(egress2_15_io_in4_3),
    .io_out4_0(egress2_15_io_out4_0),
    .io_out4_1(egress2_15_io_out4_1),
    .io_out4_2(egress2_15_io_out4_2),
    .io_out4_3(egress2_15_io_out4_3),
    .io_ctrl(egress2_15_io_ctrl)
  );
  assign io_out64_0 = egress2_0_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_1 = egress2_0_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_2 = egress2_0_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_3 = egress2_0_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_4 = egress2_1_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_5 = egress2_1_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_6 = egress2_1_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_7 = egress2_1_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_8 = egress2_2_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_9 = egress2_2_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_10 = egress2_2_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_11 = egress2_2_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_12 = egress2_3_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_13 = egress2_3_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_14 = egress2_3_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_15 = egress2_3_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_16 = egress2_4_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_17 = egress2_4_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_18 = egress2_4_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_19 = egress2_4_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_20 = egress2_5_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_21 = egress2_5_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_22 = egress2_5_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_23 = egress2_5_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_24 = egress2_6_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_25 = egress2_6_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_26 = egress2_6_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_27 = egress2_6_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_28 = egress2_7_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_29 = egress2_7_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_30 = egress2_7_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_31 = egress2_7_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_32 = egress2_8_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_33 = egress2_8_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_34 = egress2_8_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_35 = egress2_8_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_36 = egress2_9_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_37 = egress2_9_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_38 = egress2_9_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_39 = egress2_9_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_40 = egress2_10_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_41 = egress2_10_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_42 = egress2_10_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_43 = egress2_10_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_44 = egress2_11_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_45 = egress2_11_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_46 = egress2_11_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_47 = egress2_11_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_48 = egress2_12_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_49 = egress2_12_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_50 = egress2_12_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_51 = egress2_12_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_52 = egress2_13_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_53 = egress2_13_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_54 = egress2_13_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_55 = egress2_13_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_56 = egress2_14_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_57 = egress2_14_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_58 = egress2_14_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_59 = egress2_14_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_60 = egress2_15_io_out4_0[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_61 = egress2_15_io_out4_1[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_62 = egress2_15_io_out4_2[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_out64_63 = egress2_15_io_out4_3[63:0]; // @[BuildingBlock.scala 207:47]
  assign io_validout64_0 = egress2_0_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_1 = egress2_0_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_2 = egress2_0_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_3 = egress2_0_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_4 = egress2_1_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_5 = egress2_1_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_6 = egress2_1_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_7 = egress2_1_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_8 = egress2_2_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_9 = egress2_2_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_10 = egress2_2_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_11 = egress2_2_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_12 = egress2_3_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_13 = egress2_3_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_14 = egress2_3_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_15 = egress2_3_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_16 = egress2_4_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_17 = egress2_4_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_18 = egress2_4_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_19 = egress2_4_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_20 = egress2_5_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_21 = egress2_5_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_22 = egress2_5_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_23 = egress2_5_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_24 = egress2_6_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_25 = egress2_6_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_26 = egress2_6_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_27 = egress2_6_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_28 = egress2_7_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_29 = egress2_7_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_30 = egress2_7_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_31 = egress2_7_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_32 = egress2_8_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_33 = egress2_8_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_34 = egress2_8_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_35 = egress2_8_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_36 = egress2_9_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_37 = egress2_9_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_38 = egress2_9_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_39 = egress2_9_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_40 = egress2_10_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_41 = egress2_10_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_42 = egress2_10_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_43 = egress2_10_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_44 = egress2_11_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_45 = egress2_11_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_46 = egress2_11_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_47 = egress2_11_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_48 = egress2_12_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_49 = egress2_12_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_50 = egress2_12_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_51 = egress2_12_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_52 = egress2_13_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_53 = egress2_13_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_54 = egress2_13_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_55 = egress2_13_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_56 = egress2_14_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_57 = egress2_14_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_58 = egress2_14_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_59 = egress2_14_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_60 = egress2_15_io_out4_0[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_61 = egress2_15_io_out4_1[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_62 = egress2_15_io_out4_2[64]; // @[BuildingBlock.scala 208:52]
  assign io_validout64_63 = egress2_15_io_out4_3[64]; // @[BuildingBlock.scala 208:52]
  assign io_tagout_Tag = tag_Tag; // @[BuildingBlock.scala 195:13]
  assign io_tagout_RoundCnt = tag_RoundCnt; // @[BuildingBlock.scala 195:13]
  assign io_addrout = addr; // @[BuildingBlock.scala 197:14]
  assign egress2_0_clock = clock;
  assign egress2_0_io_in4_0 = {io_validin64_0,io_in64_0}; // @[Cat.scala 30:58]
  assign egress2_0_io_in4_1 = {io_validin64_1,io_in64_1}; // @[Cat.scala 30:58]
  assign egress2_0_io_in4_2 = {io_validin64_2,io_in64_2}; // @[Cat.scala 30:58]
  assign egress2_0_io_in4_3 = {io_validin64_3,io_in64_3}; // @[Cat.scala 30:58]
  assign egress2_0_io_ctrl = io_ctrl[127:120]; // @[BuildingBlock.scala 212:34]
  assign egress2_1_clock = clock;
  assign egress2_1_io_in4_0 = {io_validin64_4,io_in64_4}; // @[Cat.scala 30:58]
  assign egress2_1_io_in4_1 = {io_validin64_5,io_in64_5}; // @[Cat.scala 30:58]
  assign egress2_1_io_in4_2 = {io_validin64_6,io_in64_6}; // @[Cat.scala 30:58]
  assign egress2_1_io_in4_3 = {io_validin64_7,io_in64_7}; // @[Cat.scala 30:58]
  assign egress2_1_io_ctrl = io_ctrl[119:112]; // @[BuildingBlock.scala 212:34]
  assign egress2_2_clock = clock;
  assign egress2_2_io_in4_0 = {io_validin64_8,io_in64_8}; // @[Cat.scala 30:58]
  assign egress2_2_io_in4_1 = {io_validin64_9,io_in64_9}; // @[Cat.scala 30:58]
  assign egress2_2_io_in4_2 = {io_validin64_10,io_in64_10}; // @[Cat.scala 30:58]
  assign egress2_2_io_in4_3 = {io_validin64_11,io_in64_11}; // @[Cat.scala 30:58]
  assign egress2_2_io_ctrl = io_ctrl[111:104]; // @[BuildingBlock.scala 212:34]
  assign egress2_3_clock = clock;
  assign egress2_3_io_in4_0 = {io_validin64_12,io_in64_12}; // @[Cat.scala 30:58]
  assign egress2_3_io_in4_1 = {io_validin64_13,io_in64_13}; // @[Cat.scala 30:58]
  assign egress2_3_io_in4_2 = {io_validin64_14,io_in64_14}; // @[Cat.scala 30:58]
  assign egress2_3_io_in4_3 = {io_validin64_15,io_in64_15}; // @[Cat.scala 30:58]
  assign egress2_3_io_ctrl = io_ctrl[103:96]; // @[BuildingBlock.scala 212:34]
  assign egress2_4_clock = clock;
  assign egress2_4_io_in4_0 = {io_validin64_16,io_in64_16}; // @[Cat.scala 30:58]
  assign egress2_4_io_in4_1 = {io_validin64_17,io_in64_17}; // @[Cat.scala 30:58]
  assign egress2_4_io_in4_2 = {io_validin64_18,io_in64_18}; // @[Cat.scala 30:58]
  assign egress2_4_io_in4_3 = {io_validin64_19,io_in64_19}; // @[Cat.scala 30:58]
  assign egress2_4_io_ctrl = io_ctrl[95:88]; // @[BuildingBlock.scala 212:34]
  assign egress2_5_clock = clock;
  assign egress2_5_io_in4_0 = {io_validin64_20,io_in64_20}; // @[Cat.scala 30:58]
  assign egress2_5_io_in4_1 = {io_validin64_21,io_in64_21}; // @[Cat.scala 30:58]
  assign egress2_5_io_in4_2 = {io_validin64_22,io_in64_22}; // @[Cat.scala 30:58]
  assign egress2_5_io_in4_3 = {io_validin64_23,io_in64_23}; // @[Cat.scala 30:58]
  assign egress2_5_io_ctrl = io_ctrl[87:80]; // @[BuildingBlock.scala 212:34]
  assign egress2_6_clock = clock;
  assign egress2_6_io_in4_0 = {io_validin64_24,io_in64_24}; // @[Cat.scala 30:58]
  assign egress2_6_io_in4_1 = {io_validin64_25,io_in64_25}; // @[Cat.scala 30:58]
  assign egress2_6_io_in4_2 = {io_validin64_26,io_in64_26}; // @[Cat.scala 30:58]
  assign egress2_6_io_in4_3 = {io_validin64_27,io_in64_27}; // @[Cat.scala 30:58]
  assign egress2_6_io_ctrl = io_ctrl[79:72]; // @[BuildingBlock.scala 212:34]
  assign egress2_7_clock = clock;
  assign egress2_7_io_in4_0 = {io_validin64_28,io_in64_28}; // @[Cat.scala 30:58]
  assign egress2_7_io_in4_1 = {io_validin64_29,io_in64_29}; // @[Cat.scala 30:58]
  assign egress2_7_io_in4_2 = {io_validin64_30,io_in64_30}; // @[Cat.scala 30:58]
  assign egress2_7_io_in4_3 = {io_validin64_31,io_in64_31}; // @[Cat.scala 30:58]
  assign egress2_7_io_ctrl = io_ctrl[71:64]; // @[BuildingBlock.scala 212:34]
  assign egress2_8_clock = clock;
  assign egress2_8_io_in4_0 = {io_validin64_32,io_in64_32}; // @[Cat.scala 30:58]
  assign egress2_8_io_in4_1 = {io_validin64_33,io_in64_33}; // @[Cat.scala 30:58]
  assign egress2_8_io_in4_2 = {io_validin64_34,io_in64_34}; // @[Cat.scala 30:58]
  assign egress2_8_io_in4_3 = {io_validin64_35,io_in64_35}; // @[Cat.scala 30:58]
  assign egress2_8_io_ctrl = io_ctrl[63:56]; // @[BuildingBlock.scala 212:34]
  assign egress2_9_clock = clock;
  assign egress2_9_io_in4_0 = {io_validin64_36,io_in64_36}; // @[Cat.scala 30:58]
  assign egress2_9_io_in4_1 = {io_validin64_37,io_in64_37}; // @[Cat.scala 30:58]
  assign egress2_9_io_in4_2 = {io_validin64_38,io_in64_38}; // @[Cat.scala 30:58]
  assign egress2_9_io_in4_3 = {io_validin64_39,io_in64_39}; // @[Cat.scala 30:58]
  assign egress2_9_io_ctrl = io_ctrl[55:48]; // @[BuildingBlock.scala 212:34]
  assign egress2_10_clock = clock;
  assign egress2_10_io_in4_0 = {io_validin64_40,io_in64_40}; // @[Cat.scala 30:58]
  assign egress2_10_io_in4_1 = {io_validin64_41,io_in64_41}; // @[Cat.scala 30:58]
  assign egress2_10_io_in4_2 = {io_validin64_42,io_in64_42}; // @[Cat.scala 30:58]
  assign egress2_10_io_in4_3 = {io_validin64_43,io_in64_43}; // @[Cat.scala 30:58]
  assign egress2_10_io_ctrl = io_ctrl[47:40]; // @[BuildingBlock.scala 212:34]
  assign egress2_11_clock = clock;
  assign egress2_11_io_in4_0 = {io_validin64_44,io_in64_44}; // @[Cat.scala 30:58]
  assign egress2_11_io_in4_1 = {io_validin64_45,io_in64_45}; // @[Cat.scala 30:58]
  assign egress2_11_io_in4_2 = {io_validin64_46,io_in64_46}; // @[Cat.scala 30:58]
  assign egress2_11_io_in4_3 = {io_validin64_47,io_in64_47}; // @[Cat.scala 30:58]
  assign egress2_11_io_ctrl = io_ctrl[39:32]; // @[BuildingBlock.scala 212:34]
  assign egress2_12_clock = clock;
  assign egress2_12_io_in4_0 = {io_validin64_48,io_in64_48}; // @[Cat.scala 30:58]
  assign egress2_12_io_in4_1 = {io_validin64_49,io_in64_49}; // @[Cat.scala 30:58]
  assign egress2_12_io_in4_2 = {io_validin64_50,io_in64_50}; // @[Cat.scala 30:58]
  assign egress2_12_io_in4_3 = {io_validin64_51,io_in64_51}; // @[Cat.scala 30:58]
  assign egress2_12_io_ctrl = io_ctrl[31:24]; // @[BuildingBlock.scala 212:34]
  assign egress2_13_clock = clock;
  assign egress2_13_io_in4_0 = {io_validin64_52,io_in64_52}; // @[Cat.scala 30:58]
  assign egress2_13_io_in4_1 = {io_validin64_53,io_in64_53}; // @[Cat.scala 30:58]
  assign egress2_13_io_in4_2 = {io_validin64_54,io_in64_54}; // @[Cat.scala 30:58]
  assign egress2_13_io_in4_3 = {io_validin64_55,io_in64_55}; // @[Cat.scala 30:58]
  assign egress2_13_io_ctrl = io_ctrl[23:16]; // @[BuildingBlock.scala 212:34]
  assign egress2_14_clock = clock;
  assign egress2_14_io_in4_0 = {io_validin64_56,io_in64_56}; // @[Cat.scala 30:58]
  assign egress2_14_io_in4_1 = {io_validin64_57,io_in64_57}; // @[Cat.scala 30:58]
  assign egress2_14_io_in4_2 = {io_validin64_58,io_in64_58}; // @[Cat.scala 30:58]
  assign egress2_14_io_in4_3 = {io_validin64_59,io_in64_59}; // @[Cat.scala 30:58]
  assign egress2_14_io_ctrl = io_ctrl[15:8]; // @[BuildingBlock.scala 212:34]
  assign egress2_15_clock = clock;
  assign egress2_15_io_in4_0 = {io_validin64_60,io_in64_60}; // @[Cat.scala 30:58]
  assign egress2_15_io_in4_1 = {io_validin64_61,io_in64_61}; // @[Cat.scala 30:58]
  assign egress2_15_io_in4_2 = {io_validin64_62,io_in64_62}; // @[Cat.scala 30:58]
  assign egress2_15_io_in4_3 = {io_validin64_63,io_in64_63}; // @[Cat.scala 30:58]
  assign egress2_15_io_ctrl = io_ctrl[7:0]; // @[BuildingBlock.scala 212:34]
  always @(posedge clock) begin
    tag_Tag <= io_tagin_Tag; // @[BuildingBlock.scala 194:20]
    tag_RoundCnt <= io_tagin_RoundCnt; // @[BuildingBlock.scala 194:20]
    addr <= io_addrin; // @[BuildingBlock.scala 196:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_Tag = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  tag_RoundCnt = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  addr = _RAND_2[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BuildingBlockNew(
  input          clock,
  input          reset,
  input  [63:0]  io_d_in_0_a,
  input          io_d_in_0_valid_a,
  input  [63:0]  io_d_in_0_b,
  input  [63:0]  io_d_in_1_a,
  input          io_d_in_1_valid_a,
  input  [63:0]  io_d_in_1_b,
  input  [63:0]  io_d_in_2_a,
  input          io_d_in_2_valid_a,
  input  [63:0]  io_d_in_2_b,
  input  [63:0]  io_d_in_3_a,
  input          io_d_in_3_valid_a,
  input  [63:0]  io_d_in_3_b,
  input  [63:0]  io_d_in_4_a,
  input          io_d_in_4_valid_a,
  input  [63:0]  io_d_in_4_b,
  input  [63:0]  io_d_in_5_a,
  input          io_d_in_5_valid_a,
  input  [63:0]  io_d_in_5_b,
  input  [63:0]  io_d_in_6_a,
  input          io_d_in_6_valid_a,
  input  [63:0]  io_d_in_6_b,
  input  [63:0]  io_d_in_7_a,
  input          io_d_in_7_valid_a,
  input  [63:0]  io_d_in_7_b,
  input  [63:0]  io_d_in_8_a,
  input          io_d_in_8_valid_a,
  input  [63:0]  io_d_in_8_b,
  input  [63:0]  io_d_in_9_a,
  input          io_d_in_9_valid_a,
  input  [63:0]  io_d_in_9_b,
  input  [63:0]  io_d_in_10_a,
  input          io_d_in_10_valid_a,
  input  [63:0]  io_d_in_10_b,
  input  [63:0]  io_d_in_11_a,
  input          io_d_in_11_valid_a,
  input  [63:0]  io_d_in_11_b,
  input  [63:0]  io_d_in_12_a,
  input          io_d_in_12_valid_a,
  input  [63:0]  io_d_in_12_b,
  input  [63:0]  io_d_in_13_a,
  input          io_d_in_13_valid_a,
  input  [63:0]  io_d_in_13_b,
  input  [63:0]  io_d_in_14_a,
  input          io_d_in_14_valid_a,
  input  [63:0]  io_d_in_14_b,
  input  [63:0]  io_d_in_15_a,
  input          io_d_in_15_valid_a,
  input  [63:0]  io_d_in_15_b,
  input  [63:0]  io_d_in_16_a,
  input          io_d_in_16_valid_a,
  input  [63:0]  io_d_in_16_b,
  input  [63:0]  io_d_in_17_a,
  input          io_d_in_17_valid_a,
  input  [63:0]  io_d_in_17_b,
  input  [63:0]  io_d_in_18_a,
  input          io_d_in_18_valid_a,
  input  [63:0]  io_d_in_18_b,
  input  [63:0]  io_d_in_19_a,
  input          io_d_in_19_valid_a,
  input  [63:0]  io_d_in_19_b,
  input  [63:0]  io_d_in_20_a,
  input          io_d_in_20_valid_a,
  input  [63:0]  io_d_in_20_b,
  input  [63:0]  io_d_in_21_a,
  input          io_d_in_21_valid_a,
  input  [63:0]  io_d_in_21_b,
  input  [63:0]  io_d_in_22_a,
  input          io_d_in_22_valid_a,
  input  [63:0]  io_d_in_22_b,
  input  [63:0]  io_d_in_23_a,
  input          io_d_in_23_valid_a,
  input  [63:0]  io_d_in_23_b,
  input  [63:0]  io_d_in_24_a,
  input          io_d_in_24_valid_a,
  input  [63:0]  io_d_in_24_b,
  input  [63:0]  io_d_in_25_a,
  input          io_d_in_25_valid_a,
  input  [63:0]  io_d_in_25_b,
  input  [63:0]  io_d_in_26_a,
  input          io_d_in_26_valid_a,
  input  [63:0]  io_d_in_26_b,
  input  [63:0]  io_d_in_27_a,
  input          io_d_in_27_valid_a,
  input  [63:0]  io_d_in_27_b,
  input  [63:0]  io_d_in_28_a,
  input          io_d_in_28_valid_a,
  input  [63:0]  io_d_in_28_b,
  input  [63:0]  io_d_in_29_a,
  input          io_d_in_29_valid_a,
  input  [63:0]  io_d_in_29_b,
  input  [63:0]  io_d_in_30_a,
  input          io_d_in_30_valid_a,
  input  [63:0]  io_d_in_30_b,
  input  [63:0]  io_d_in_31_a,
  input          io_d_in_31_valid_a,
  input  [63:0]  io_d_in_31_b,
  output [63:0]  io_d_out_0_a,
  output         io_d_out_0_valid_a,
  output [63:0]  io_d_out_0_b,
  output         io_d_out_0_valid_b,
  output [63:0]  io_d_out_1_a,
  output         io_d_out_1_valid_a,
  output [63:0]  io_d_out_1_b,
  output         io_d_out_1_valid_b,
  output [63:0]  io_d_out_2_a,
  output         io_d_out_2_valid_a,
  output [63:0]  io_d_out_2_b,
  output         io_d_out_2_valid_b,
  output [63:0]  io_d_out_3_a,
  output         io_d_out_3_valid_a,
  output [63:0]  io_d_out_3_b,
  output         io_d_out_3_valid_b,
  output [63:0]  io_d_out_4_a,
  output         io_d_out_4_valid_a,
  output [63:0]  io_d_out_4_b,
  output         io_d_out_4_valid_b,
  output [63:0]  io_d_out_5_a,
  output         io_d_out_5_valid_a,
  output [63:0]  io_d_out_5_b,
  output         io_d_out_5_valid_b,
  output [63:0]  io_d_out_6_a,
  output         io_d_out_6_valid_a,
  output [63:0]  io_d_out_6_b,
  output         io_d_out_6_valid_b,
  output [63:0]  io_d_out_7_a,
  output         io_d_out_7_valid_a,
  output [63:0]  io_d_out_7_b,
  output         io_d_out_7_valid_b,
  output [63:0]  io_d_out_8_a,
  output         io_d_out_8_valid_a,
  output [63:0]  io_d_out_8_b,
  output         io_d_out_8_valid_b,
  output [63:0]  io_d_out_9_a,
  output         io_d_out_9_valid_a,
  output [63:0]  io_d_out_9_b,
  output         io_d_out_9_valid_b,
  output [63:0]  io_d_out_10_a,
  output         io_d_out_10_valid_a,
  output [63:0]  io_d_out_10_b,
  output         io_d_out_10_valid_b,
  output [63:0]  io_d_out_11_a,
  output         io_d_out_11_valid_a,
  output [63:0]  io_d_out_11_b,
  output         io_d_out_11_valid_b,
  output [63:0]  io_d_out_12_a,
  output         io_d_out_12_valid_a,
  output [63:0]  io_d_out_12_b,
  output         io_d_out_12_valid_b,
  output [63:0]  io_d_out_13_a,
  output         io_d_out_13_valid_a,
  output [63:0]  io_d_out_13_b,
  output         io_d_out_13_valid_b,
  output [63:0]  io_d_out_14_a,
  output         io_d_out_14_valid_a,
  output [63:0]  io_d_out_14_b,
  output         io_d_out_14_valid_b,
  output [63:0]  io_d_out_15_a,
  output         io_d_out_15_valid_a,
  output [63:0]  io_d_out_15_b,
  output         io_d_out_15_valid_b,
  output [63:0]  io_d_out_16_a,
  output         io_d_out_16_valid_a,
  output [63:0]  io_d_out_16_b,
  output         io_d_out_16_valid_b,
  output [63:0]  io_d_out_17_a,
  output         io_d_out_17_valid_a,
  output [63:0]  io_d_out_17_b,
  output         io_d_out_17_valid_b,
  output [63:0]  io_d_out_18_a,
  output         io_d_out_18_valid_a,
  output [63:0]  io_d_out_18_b,
  output         io_d_out_18_valid_b,
  output [63:0]  io_d_out_19_a,
  output         io_d_out_19_valid_a,
  output [63:0]  io_d_out_19_b,
  output         io_d_out_19_valid_b,
  output [63:0]  io_d_out_20_a,
  output         io_d_out_20_valid_a,
  output [63:0]  io_d_out_20_b,
  output         io_d_out_20_valid_b,
  output [63:0]  io_d_out_21_a,
  output         io_d_out_21_valid_a,
  output [63:0]  io_d_out_21_b,
  output         io_d_out_21_valid_b,
  output [63:0]  io_d_out_22_a,
  output         io_d_out_22_valid_a,
  output [63:0]  io_d_out_22_b,
  output         io_d_out_22_valid_b,
  output [63:0]  io_d_out_23_a,
  output         io_d_out_23_valid_a,
  output [63:0]  io_d_out_23_b,
  output         io_d_out_23_valid_b,
  output [63:0]  io_d_out_24_a,
  output         io_d_out_24_valid_a,
  output [63:0]  io_d_out_24_b,
  output         io_d_out_24_valid_b,
  output [63:0]  io_d_out_25_a,
  output         io_d_out_25_valid_a,
  output [63:0]  io_d_out_25_b,
  output         io_d_out_25_valid_b,
  output [63:0]  io_d_out_26_a,
  output         io_d_out_26_valid_a,
  output [63:0]  io_d_out_26_b,
  output         io_d_out_26_valid_b,
  output [63:0]  io_d_out_27_a,
  output         io_d_out_27_valid_a,
  output [63:0]  io_d_out_27_b,
  output         io_d_out_27_valid_b,
  output [63:0]  io_d_out_28_a,
  output         io_d_out_28_valid_a,
  output [63:0]  io_d_out_28_b,
  output         io_d_out_28_valid_b,
  output [63:0]  io_d_out_29_a,
  output         io_d_out_29_valid_a,
  output [63:0]  io_d_out_29_b,
  output         io_d_out_29_valid_b,
  output [63:0]  io_d_out_30_a,
  output         io_d_out_30_valid_a,
  output [63:0]  io_d_out_30_b,
  output         io_d_out_30_valid_b,
  output [63:0]  io_d_out_31_a,
  output         io_d_out_31_valid_a,
  output [63:0]  io_d_out_31_b,
  output         io_d_out_31_valid_b,
  input          io_wr_en_mem1,
  input          io_wr_en_mem2,
  input          io_wr_en_mem3,
  input          io_wr_en_mem4,
  input          io_wr_en_mem5,
  input          io_wr_en_mem6,
  input  [287:0] io_wr_instr_mem1,
  input  [127:0] io_wr_instr_mem2,
  input  [127:0] io_wr_instr_mem3,
  input  [127:0] io_wr_instr_mem4,
  input  [127:0] io_wr_instr_mem5,
  input  [127:0] io_wr_instr_mem6,
  input  [7:0]   io_PC1_in,
  output [7:0]   io_PC6_out,
  input  [7:0]   io_Addr_in,
  output [7:0]   io_Addr_out,
  input  [1:0]   io_Tag_in_Tag,
  input  [2:0]   io_Tag_in_RoundCnt,
  output [1:0]   io_Tag_out_Tag,
  output [2:0]   io_Tag_out_RoundCnt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [287:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [127:0] _RAND_14;
  reg [127:0] _RAND_15;
  reg [127:0] _RAND_16;
  reg [127:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] Mem1_R0_addr; // @[BuildingBlockNew.scala 34:25]
  wire  Mem1_R0_clk; // @[BuildingBlockNew.scala 34:25]
  wire [287:0] Mem1_R0_data; // @[BuildingBlockNew.scala 34:25]
  wire [7:0] Mem1_W0_addr; // @[BuildingBlockNew.scala 34:25]
  wire  Mem1_W0_en; // @[BuildingBlockNew.scala 34:25]
  wire  Mem1_W0_clk; // @[BuildingBlockNew.scala 34:25]
  wire [287:0] Mem1_W0_data; // @[BuildingBlockNew.scala 34:25]
  wire [7:0] Mem2_R0_addr; // @[BuildingBlockNew.scala 35:25]
  wire  Mem2_R0_clk; // @[BuildingBlockNew.scala 35:25]
  wire [127:0] Mem2_R0_data; // @[BuildingBlockNew.scala 35:25]
  wire [7:0] Mem2_W0_addr; // @[BuildingBlockNew.scala 35:25]
  wire  Mem2_W0_en; // @[BuildingBlockNew.scala 35:25]
  wire  Mem2_W0_clk; // @[BuildingBlockNew.scala 35:25]
  wire [127:0] Mem2_W0_data; // @[BuildingBlockNew.scala 35:25]
  wire [7:0] Mem3_R0_addr; // @[BuildingBlockNew.scala 36:25]
  wire  Mem3_R0_clk; // @[BuildingBlockNew.scala 36:25]
  wire [127:0] Mem3_R0_data; // @[BuildingBlockNew.scala 36:25]
  wire [7:0] Mem3_W0_addr; // @[BuildingBlockNew.scala 36:25]
  wire  Mem3_W0_en; // @[BuildingBlockNew.scala 36:25]
  wire  Mem3_W0_clk; // @[BuildingBlockNew.scala 36:25]
  wire [127:0] Mem3_W0_data; // @[BuildingBlockNew.scala 36:25]
  wire [7:0] Mem4_R0_addr; // @[BuildingBlockNew.scala 37:25]
  wire  Mem4_R0_clk; // @[BuildingBlockNew.scala 37:25]
  wire [127:0] Mem4_R0_data; // @[BuildingBlockNew.scala 37:25]
  wire [7:0] Mem4_W0_addr; // @[BuildingBlockNew.scala 37:25]
  wire  Mem4_W0_en; // @[BuildingBlockNew.scala 37:25]
  wire  Mem4_W0_clk; // @[BuildingBlockNew.scala 37:25]
  wire [127:0] Mem4_W0_data; // @[BuildingBlockNew.scala 37:25]
  wire [7:0] Mem5_R0_addr; // @[BuildingBlockNew.scala 38:25]
  wire  Mem5_R0_clk; // @[BuildingBlockNew.scala 38:25]
  wire [127:0] Mem5_R0_data; // @[BuildingBlockNew.scala 38:25]
  wire [7:0] Mem5_W0_addr; // @[BuildingBlockNew.scala 38:25]
  wire  Mem5_W0_en; // @[BuildingBlockNew.scala 38:25]
  wire  Mem5_W0_clk; // @[BuildingBlockNew.scala 38:25]
  wire [127:0] Mem5_W0_data; // @[BuildingBlockNew.scala 38:25]
  wire [7:0] Mem6_R0_addr; // @[BuildingBlockNew.scala 39:25]
  wire  Mem6_R0_clk; // @[BuildingBlockNew.scala 39:25]
  wire [127:0] Mem6_R0_data; // @[BuildingBlockNew.scala 39:25]
  wire [7:0] Mem6_W0_addr; // @[BuildingBlockNew.scala 39:25]
  wire  Mem6_W0_en; // @[BuildingBlockNew.scala 39:25]
  wire  Mem6_W0_clk; // @[BuildingBlockNew.scala 39:25]
  wire [127:0] Mem6_W0_data; // @[BuildingBlockNew.scala 39:25]
  wire  peCol_clock; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_reset; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_0_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_0_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_0_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_1_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_1_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_1_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_2_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_2_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_2_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_3_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_3_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_3_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_4_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_4_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_4_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_5_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_5_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_5_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_6_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_6_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_6_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_7_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_7_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_7_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_8_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_8_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_8_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_9_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_9_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_9_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_10_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_10_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_10_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_11_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_11_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_11_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_12_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_12_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_12_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_13_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_13_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_13_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_14_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_14_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_14_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_15_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_15_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_15_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_16_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_16_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_16_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_17_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_17_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_17_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_18_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_18_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_18_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_19_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_19_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_19_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_20_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_20_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_20_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_21_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_21_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_21_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_22_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_22_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_22_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_23_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_23_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_23_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_24_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_24_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_24_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_25_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_25_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_25_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_26_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_26_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_26_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_27_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_27_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_27_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_28_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_28_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_28_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_29_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_29_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_29_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_30_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_30_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_30_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_31_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_31_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_in_31_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_0_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_0_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_0_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_1_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_1_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_1_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_2_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_2_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_2_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_3_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_3_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_3_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_4_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_4_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_4_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_5_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_5_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_5_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_6_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_6_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_6_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_7_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_7_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_7_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_8_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_8_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_8_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_9_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_9_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_9_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_10_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_10_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_10_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_11_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_11_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_11_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_12_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_12_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_12_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_13_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_13_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_13_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_14_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_14_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_14_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_15_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_15_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_15_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_16_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_16_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_16_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_17_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_17_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_17_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_18_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_18_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_18_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_19_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_19_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_19_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_20_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_20_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_20_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_21_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_21_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_21_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_22_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_22_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_22_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_23_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_23_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_23_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_24_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_24_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_24_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_25_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_25_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_25_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_26_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_26_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_26_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_27_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_27_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_27_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_28_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_28_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_28_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_29_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_29_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_29_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_30_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_30_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_30_b; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_31_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_31_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [63:0] peCol_io_d_out_31_b; // @[BuildingBlockNew.scala 83:21]
  wire [1:0] peCol_io_tagin_Tag; // @[BuildingBlockNew.scala 83:21]
  wire [2:0] peCol_io_tagin_RoundCnt; // @[BuildingBlockNew.scala 83:21]
  wire [7:0] peCol_io_addrin; // @[BuildingBlockNew.scala 83:21]
  wire [1:0] peCol_io_tagout_Tag; // @[BuildingBlockNew.scala 83:21]
  wire [2:0] peCol_io_tagout_RoundCnt; // @[BuildingBlockNew.scala 83:21]
  wire [7:0] peCol_io_addrout; // @[BuildingBlockNew.scala 83:21]
  wire [287:0] peCol_io_instr; // @[BuildingBlockNew.scala 83:21]
  wire  ingress1_clock; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_0; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_1; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_2; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_3; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_4; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_5; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_6; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_7; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_8; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_9; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_10; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_11; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_12; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_13; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_14; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_15; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_16; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_17; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_18; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_19; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_20; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_21; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_22; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_23; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_24; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_25; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_26; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_27; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_28; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_29; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_30; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_31; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_32; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_33; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_34; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_35; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_36; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_37; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_38; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_39; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_40; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_41; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_42; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_43; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_44; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_45; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_46; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_47; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_48; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_49; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_50; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_51; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_52; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_53; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_54; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_55; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_56; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_57; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_58; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_59; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_60; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_61; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_62; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_in64_63; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_0; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_2; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_4; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_6; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_8; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_10; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_12; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_14; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_16; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_18; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_20; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_22; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_24; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_26; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_28; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_30; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_32; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_34; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_36; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_38; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_40; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_42; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_44; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_46; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_48; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_50; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_52; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_54; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_56; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_58; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_60; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_62; // @[BuildingBlockNew.scala 84:24]
  wire [1:0] ingress1_io_tagin_Tag; // @[BuildingBlockNew.scala 84:24]
  wire [2:0] ingress1_io_tagin_RoundCnt; // @[BuildingBlockNew.scala 84:24]
  wire [7:0] ingress1_io_addrin; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_0; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_1; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_2; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_3; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_4; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_5; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_6; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_7; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_8; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_9; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_10; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_11; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_12; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_13; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_14; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_15; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_16; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_17; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_18; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_19; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_20; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_21; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_22; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_23; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_24; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_25; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_26; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_27; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_28; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_29; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_30; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_31; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_32; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_33; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_34; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_35; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_36; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_37; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_38; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_39; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_40; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_41; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_42; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_43; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_44; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_45; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_46; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_47; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_48; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_49; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_50; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_51; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_52; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_53; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_54; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_55; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_56; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_57; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_58; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_59; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_60; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_61; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_62; // @[BuildingBlockNew.scala 84:24]
  wire [63:0] ingress1_io_out64_63; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_0; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_1; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_2; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_3; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_4; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_5; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_6; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_7; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_8; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_9; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_10; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_11; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_12; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_13; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_14; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_15; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_16; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_17; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_18; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_19; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_20; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_21; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_22; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_23; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_24; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_25; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_26; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_27; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_28; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_29; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_30; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_31; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_32; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_33; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_34; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_35; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_36; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_37; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_38; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_39; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_40; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_41; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_42; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_43; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_44; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_45; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_46; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_47; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_48; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_49; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_50; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_51; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_52; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_53; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_54; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_55; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_56; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_57; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_58; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_59; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_60; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_61; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_62; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_63; // @[BuildingBlockNew.scala 84:24]
  wire [1:0] ingress1_io_tagout_Tag; // @[BuildingBlockNew.scala 84:24]
  wire [2:0] ingress1_io_tagout_RoundCnt; // @[BuildingBlockNew.scala 84:24]
  wire [7:0] ingress1_io_addrout; // @[BuildingBlockNew.scala 84:24]
  wire [127:0] ingress1_io_ctrl; // @[BuildingBlockNew.scala 84:24]
  wire  ingress2_clock; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_0; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_1; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_2; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_3; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_4; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_5; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_6; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_7; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_8; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_9; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_10; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_11; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_12; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_13; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_14; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_15; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_16; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_17; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_18; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_19; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_20; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_21; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_22; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_23; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_24; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_25; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_26; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_27; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_28; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_29; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_30; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_31; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_32; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_33; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_34; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_35; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_36; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_37; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_38; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_39; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_40; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_41; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_42; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_43; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_44; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_45; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_46; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_47; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_48; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_49; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_50; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_51; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_52; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_53; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_54; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_55; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_56; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_57; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_58; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_59; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_60; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_61; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_62; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_in64_63; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_0; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_1; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_2; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_3; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_4; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_5; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_6; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_7; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_8; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_9; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_10; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_11; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_12; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_13; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_14; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_15; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_16; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_17; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_18; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_19; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_20; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_21; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_22; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_23; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_24; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_25; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_26; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_27; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_28; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_29; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_30; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_31; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_32; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_33; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_34; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_35; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_36; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_37; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_38; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_39; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_40; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_41; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_42; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_43; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_44; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_45; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_46; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_47; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_48; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_49; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_50; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_51; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_52; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_53; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_54; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_55; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_56; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_57; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_58; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_59; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_60; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_61; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_62; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_63; // @[BuildingBlockNew.scala 85:24]
  wire [1:0] ingress2_io_tagin_Tag; // @[BuildingBlockNew.scala 85:24]
  wire [2:0] ingress2_io_tagin_RoundCnt; // @[BuildingBlockNew.scala 85:24]
  wire [7:0] ingress2_io_addrin; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_0; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_1; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_2; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_3; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_4; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_5; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_6; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_7; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_8; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_9; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_10; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_11; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_12; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_13; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_14; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_15; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_16; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_17; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_18; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_19; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_20; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_21; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_22; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_23; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_24; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_25; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_26; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_27; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_28; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_29; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_30; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_31; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_32; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_33; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_34; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_35; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_36; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_37; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_38; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_39; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_40; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_41; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_42; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_43; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_44; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_45; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_46; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_47; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_48; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_49; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_50; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_51; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_52; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_53; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_54; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_55; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_56; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_57; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_58; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_59; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_60; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_61; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_62; // @[BuildingBlockNew.scala 85:24]
  wire [63:0] ingress2_io_out64_63; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_0; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_1; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_2; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_3; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_4; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_5; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_6; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_7; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_8; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_9; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_10; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_11; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_12; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_13; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_14; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_15; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_16; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_17; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_18; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_19; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_20; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_21; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_22; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_23; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_24; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_25; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_26; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_27; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_28; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_29; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_30; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_31; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_32; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_33; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_34; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_35; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_36; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_37; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_38; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_39; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_40; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_41; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_42; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_43; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_44; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_45; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_46; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_47; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_48; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_49; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_50; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_51; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_52; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_53; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_54; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_55; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_56; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_57; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_58; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_59; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_60; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_61; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_62; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_63; // @[BuildingBlockNew.scala 85:24]
  wire [1:0] ingress2_io_tagout_Tag; // @[BuildingBlockNew.scala 85:24]
  wire [2:0] ingress2_io_tagout_RoundCnt; // @[BuildingBlockNew.scala 85:24]
  wire [7:0] ingress2_io_addrout; // @[BuildingBlockNew.scala 85:24]
  wire [127:0] ingress2_io_ctrl; // @[BuildingBlockNew.scala 85:24]
  wire  middle_clock; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_0; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_1; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_2; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_3; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_4; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_5; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_6; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_7; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_8; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_9; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_10; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_11; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_12; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_13; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_14; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_15; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_16; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_17; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_18; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_19; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_20; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_21; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_22; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_23; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_24; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_25; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_26; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_27; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_28; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_29; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_30; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_31; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_32; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_33; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_34; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_35; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_36; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_37; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_38; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_39; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_40; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_41; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_42; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_43; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_44; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_45; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_46; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_47; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_48; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_49; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_50; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_51; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_52; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_53; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_54; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_55; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_56; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_57; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_58; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_59; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_60; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_61; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_62; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_in64_63; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_0; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_1; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_2; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_3; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_4; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_5; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_6; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_7; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_8; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_9; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_10; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_11; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_12; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_13; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_14; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_15; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_16; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_17; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_18; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_19; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_20; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_21; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_22; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_23; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_24; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_25; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_26; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_27; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_28; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_29; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_30; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_31; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_32; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_33; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_34; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_35; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_36; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_37; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_38; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_39; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_40; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_41; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_42; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_43; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_44; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_45; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_46; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_47; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_48; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_49; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_50; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_51; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_52; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_53; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_54; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_55; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_56; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_57; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_58; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_59; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_60; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_61; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_62; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_63; // @[BuildingBlockNew.scala 86:22]
  wire [1:0] middle_io_tagin_Tag; // @[BuildingBlockNew.scala 86:22]
  wire [2:0] middle_io_tagin_RoundCnt; // @[BuildingBlockNew.scala 86:22]
  wire [7:0] middle_io_addrin; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_0; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_1; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_2; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_3; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_4; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_5; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_6; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_7; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_8; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_9; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_10; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_11; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_12; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_13; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_14; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_15; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_16; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_17; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_18; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_19; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_20; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_21; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_22; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_23; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_24; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_25; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_26; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_27; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_28; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_29; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_30; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_31; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_32; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_33; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_34; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_35; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_36; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_37; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_38; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_39; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_40; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_41; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_42; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_43; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_44; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_45; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_46; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_47; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_48; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_49; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_50; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_51; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_52; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_53; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_54; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_55; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_56; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_57; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_58; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_59; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_60; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_61; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_62; // @[BuildingBlockNew.scala 86:22]
  wire [63:0] middle_io_out64_63; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_0; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_1; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_2; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_3; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_4; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_5; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_6; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_7; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_8; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_9; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_10; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_11; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_12; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_13; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_14; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_15; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_16; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_17; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_18; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_19; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_20; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_21; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_22; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_23; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_24; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_25; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_26; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_27; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_28; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_29; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_30; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_31; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_32; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_33; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_34; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_35; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_36; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_37; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_38; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_39; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_40; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_41; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_42; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_43; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_44; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_45; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_46; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_47; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_48; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_49; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_50; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_51; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_52; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_53; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_54; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_55; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_56; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_57; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_58; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_59; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_60; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_61; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_62; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_63; // @[BuildingBlockNew.scala 86:22]
  wire [1:0] middle_io_tagout_Tag; // @[BuildingBlockNew.scala 86:22]
  wire [2:0] middle_io_tagout_RoundCnt; // @[BuildingBlockNew.scala 86:22]
  wire [7:0] middle_io_addrout; // @[BuildingBlockNew.scala 86:22]
  wire [127:0] middle_io_ctrl; // @[BuildingBlockNew.scala 86:22]
  wire  egress1_clock; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_0; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_1; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_2; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_3; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_4; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_5; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_6; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_7; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_8; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_9; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_10; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_11; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_12; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_13; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_14; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_15; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_16; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_17; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_18; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_19; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_20; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_21; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_22; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_23; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_24; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_25; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_26; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_27; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_28; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_29; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_30; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_31; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_32; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_33; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_34; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_35; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_36; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_37; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_38; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_39; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_40; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_41; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_42; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_43; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_44; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_45; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_46; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_47; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_48; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_49; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_50; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_51; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_52; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_53; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_54; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_55; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_56; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_57; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_58; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_59; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_60; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_61; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_62; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_in64_63; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_0; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_1; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_2; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_3; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_4; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_5; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_6; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_7; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_8; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_9; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_10; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_11; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_12; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_13; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_14; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_15; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_16; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_17; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_18; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_19; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_20; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_21; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_22; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_23; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_24; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_25; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_26; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_27; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_28; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_29; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_30; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_31; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_32; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_33; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_34; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_35; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_36; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_37; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_38; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_39; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_40; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_41; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_42; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_43; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_44; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_45; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_46; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_47; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_48; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_49; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_50; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_51; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_52; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_53; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_54; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_55; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_56; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_57; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_58; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_59; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_60; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_61; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_62; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_63; // @[BuildingBlockNew.scala 87:23]
  wire [1:0] egress1_io_tagin_Tag; // @[BuildingBlockNew.scala 87:23]
  wire [2:0] egress1_io_tagin_RoundCnt; // @[BuildingBlockNew.scala 87:23]
  wire [7:0] egress1_io_addrin; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_0; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_1; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_2; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_3; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_4; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_5; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_6; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_7; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_8; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_9; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_10; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_11; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_12; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_13; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_14; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_15; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_16; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_17; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_18; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_19; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_20; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_21; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_22; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_23; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_24; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_25; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_26; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_27; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_28; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_29; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_30; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_31; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_32; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_33; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_34; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_35; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_36; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_37; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_38; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_39; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_40; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_41; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_42; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_43; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_44; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_45; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_46; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_47; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_48; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_49; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_50; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_51; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_52; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_53; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_54; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_55; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_56; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_57; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_58; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_59; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_60; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_61; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_62; // @[BuildingBlockNew.scala 87:23]
  wire [63:0] egress1_io_out64_63; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_0; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_1; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_2; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_3; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_4; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_5; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_6; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_7; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_8; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_9; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_10; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_11; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_12; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_13; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_14; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_15; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_16; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_17; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_18; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_19; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_20; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_21; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_22; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_23; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_24; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_25; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_26; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_27; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_28; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_29; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_30; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_31; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_32; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_33; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_34; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_35; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_36; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_37; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_38; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_39; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_40; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_41; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_42; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_43; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_44; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_45; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_46; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_47; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_48; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_49; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_50; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_51; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_52; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_53; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_54; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_55; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_56; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_57; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_58; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_59; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_60; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_61; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_62; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_63; // @[BuildingBlockNew.scala 87:23]
  wire [1:0] egress1_io_tagout_Tag; // @[BuildingBlockNew.scala 87:23]
  wire [2:0] egress1_io_tagout_RoundCnt; // @[BuildingBlockNew.scala 87:23]
  wire [7:0] egress1_io_addrout; // @[BuildingBlockNew.scala 87:23]
  wire [127:0] egress1_io_ctrl; // @[BuildingBlockNew.scala 87:23]
  wire  egress2_clock; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_0; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_1; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_2; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_3; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_4; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_5; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_6; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_7; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_8; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_9; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_10; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_11; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_12; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_13; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_14; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_15; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_16; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_17; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_18; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_19; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_20; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_21; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_22; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_23; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_24; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_25; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_26; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_27; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_28; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_29; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_30; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_31; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_32; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_33; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_34; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_35; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_36; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_37; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_38; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_39; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_40; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_41; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_42; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_43; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_44; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_45; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_46; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_47; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_48; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_49; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_50; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_51; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_52; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_53; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_54; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_55; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_56; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_57; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_58; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_59; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_60; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_61; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_62; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_in64_63; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_0; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_1; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_2; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_3; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_4; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_5; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_6; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_7; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_8; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_9; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_10; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_11; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_12; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_13; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_14; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_15; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_16; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_17; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_18; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_19; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_20; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_21; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_22; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_23; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_24; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_25; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_26; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_27; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_28; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_29; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_30; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_31; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_32; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_33; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_34; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_35; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_36; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_37; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_38; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_39; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_40; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_41; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_42; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_43; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_44; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_45; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_46; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_47; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_48; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_49; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_50; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_51; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_52; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_53; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_54; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_55; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_56; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_57; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_58; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_59; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_60; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_61; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_62; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_63; // @[BuildingBlockNew.scala 88:23]
  wire [1:0] egress2_io_tagin_Tag; // @[BuildingBlockNew.scala 88:23]
  wire [2:0] egress2_io_tagin_RoundCnt; // @[BuildingBlockNew.scala 88:23]
  wire [7:0] egress2_io_addrin; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_0; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_1; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_2; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_3; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_4; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_5; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_6; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_7; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_8; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_9; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_10; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_11; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_12; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_13; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_14; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_15; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_16; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_17; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_18; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_19; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_20; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_21; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_22; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_23; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_24; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_25; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_26; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_27; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_28; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_29; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_30; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_31; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_32; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_33; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_34; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_35; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_36; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_37; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_38; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_39; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_40; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_41; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_42; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_43; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_44; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_45; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_46; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_47; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_48; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_49; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_50; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_51; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_52; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_53; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_54; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_55; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_56; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_57; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_58; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_59; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_60; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_61; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_62; // @[BuildingBlockNew.scala 88:23]
  wire [63:0] egress2_io_out64_63; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_0; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_1; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_2; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_3; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_4; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_5; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_6; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_7; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_8; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_9; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_10; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_11; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_12; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_13; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_14; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_15; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_16; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_17; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_18; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_19; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_20; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_21; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_22; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_23; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_24; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_25; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_26; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_27; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_28; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_29; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_30; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_31; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_32; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_33; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_34; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_35; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_36; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_37; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_38; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_39; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_40; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_41; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_42; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_43; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_44; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_45; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_46; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_47; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_48; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_49; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_50; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_51; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_52; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_53; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_54; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_55; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_56; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_57; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_58; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_59; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_60; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_61; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_62; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_63; // @[BuildingBlockNew.scala 88:23]
  wire [1:0] egress2_io_tagout_Tag; // @[BuildingBlockNew.scala 88:23]
  wire [2:0] egress2_io_tagout_RoundCnt; // @[BuildingBlockNew.scala 88:23]
  wire [7:0] egress2_io_addrout; // @[BuildingBlockNew.scala 88:23]
  wire [127:0] egress2_io_ctrl; // @[BuildingBlockNew.scala 88:23]
  reg [7:0] PC1; // @[BuildingBlockNew.scala 40:20]
  reg [7:0] PC2; // @[BuildingBlockNew.scala 41:20]
  reg [7:0] PC3; // @[BuildingBlockNew.scala 42:20]
  reg [7:0] PC4; // @[BuildingBlockNew.scala 43:20]
  reg [7:0] PC5; // @[BuildingBlockNew.scala 44:20]
  reg [7:0] PC6; // @[BuildingBlockNew.scala 45:20]
  reg [7:0] wrAddr1; // @[BuildingBlockNew.scala 46:24]
  reg [7:0] wrAddr2; // @[BuildingBlockNew.scala 47:24]
  reg [7:0] wrAddr3; // @[BuildingBlockNew.scala 48:24]
  reg [7:0] wrAddr4; // @[BuildingBlockNew.scala 49:24]
  reg [7:0] wrAddr5; // @[BuildingBlockNew.scala 50:24]
  reg [7:0] wrAddr6; // @[BuildingBlockNew.scala 51:24]
  reg [287:0] instr1; // @[BuildingBlockNew.scala 53:21]
  reg [127:0] instr2; // @[BuildingBlockNew.scala 54:21]
  reg [127:0] instr3; // @[BuildingBlockNew.scala 55:21]
  reg [127:0] instr4; // @[BuildingBlockNew.scala 56:21]
  reg [127:0] instr5; // @[BuildingBlockNew.scala 57:21]
  reg [127:0] instr6; // @[BuildingBlockNew.scala 58:21]
  wire [7:0] _wrAddr1_T_1 = wrAddr1 + 8'h1; // @[BuildingBlockNew.scala 226:24]
  wire [7:0] _wrAddr2_T_1 = wrAddr2 + 8'h1; // @[BuildingBlockNew.scala 235:24]
  wire [7:0] _wrAddr3_T_1 = wrAddr3 + 8'h1; // @[BuildingBlockNew.scala 244:24]
  wire [7:0] _wrAddr4_T_1 = wrAddr4 + 8'h1; // @[BuildingBlockNew.scala 253:24]
  wire [7:0] _wrAddr5_T_1 = wrAddr5 + 8'h1; // @[BuildingBlockNew.scala 262:24]
  wire [7:0] _wrAddr6_T_1 = wrAddr6 + 8'h1; // @[BuildingBlockNew.scala 271:24]
    sram_288_256_scn4m_subm Mem1 ( // @[BuildingBlockNew.scala 34:25]
      //.R0_addr(Mem1_R0_addr),
      //.R0_clk(Mem1_R0_clk),
      //.R0_data(Mem1_R0_data),
      //.W0_addr(Mem1_W0_addr),
      //.W0_en(Mem1_W0_en),
      //.W0_clk(Mem1_W0_clk),
      //.W0_data(Mem1_W0_data)

      //W
      .clk0(Mem1_W0_clk),
      .csb0(~Mem1_W0_en),
      .addr0(Mem1_W0_addr),
      .din0(Mem1_W0_data),
      //R
      .clk1(Mem1_R0_clk),
      .csb1(1'b0),
      .addr1(Mem1_R0_addr),
      .dout1(Mem1_R0_data)

    );
    sram_128_256_scn4m_subm Mem2 ( // @[BuildingBlockNew.scala 35:25]
      //.R0_addr(Mem2_R0_addr),
      //.R0_clk(Mem2_R0_clk),
      //.R0_data(Mem2_R0_data),
      //.W0_addr(Mem2_W0_addr),
      //.W0_en(Mem2_W0_en),
      //.W0_clk(Mem2_W0_clk),
      //.W0_data(Mem2_W0_data)

      //W
      .clk0(Mem2_W0_clk),
      .csb0(~Mem2_W0_en),
      .addr0(Mem2_W0_addr),
      .din0(Mem2_W0_data),
      //R
      .clk1(Mem2_R0_clk),
      .csb1(1'b0),
      .addr1(Mem2_R0_addr),
      .dout1(Mem2_R0_data)
    );
    sram_128_256_scn4m_subm Mem3 ( // @[BuildingBlockNew.scala 36:25]
      // .R0_addr(Mem3_R0_addr),
      // .R0_clk(Mem3_R0_clk),
      // .R0_data(Mem3_R0_data),
      // .W0_addr(Mem3_W0_addr),
      // .W0_en(Mem3_W0_en),
      // .W0_clk(Mem3_W0_clk),
      // .W0_data(Mem3_W0_data)

      //W
      .clk0(Mem3_W0_clk),
      .csb0(~Mem3_W0_en),
      .addr0(Mem3_W0_addr),
      .din0(Mem3_W0_data),
      //R
      .clk1(Mem3_R0_clk),
      .csb1(1'b0),
      .addr1(Mem3_R0_addr),
      .dout1(Mem3_R0_data)
    );
    sram_128_256_scn4m_subm Mem4 ( // @[BuildingBlockNew.scala 37:25]
      // .R0_addr(Mem4_R0_addr),
      // .R0_clk(Mem4_R0_clk),
      // .R0_data(Mem4_R0_data),
      // .W0_addr(Mem4_W0_addr),
      // .W0_en(Mem4_W0_en),
      // .W0_clk(Mem4_W0_clk),
      // .W0_data(Mem4_W0_data)

      //W
      .clk0(Mem4_W0_clk),
      .csb0(~Mem4_W0_en),
      .addr0(Mem4_W0_addr),
      .din0(Mem4_W0_data),
      //R
      .clk1(Mem4_R0_clk),
      .csb1(1'b0),
      .addr1(Mem4_R0_addr),
      .dout1(Mem4_R0_data)
    );
    sram_128_256_scn4m_subm Mem5 ( // @[BuildingBlockNew.scala 38:25]
      // .R0_addr(Mem5_R0_addr),
      // .R0_clk(Mem5_R0_clk),
      // .R0_data(Mem5_R0_data),
      // .W0_addr(Mem5_W0_addr),
      // .W0_en(Mem5_W0_en),
      // .W0_clk(Mem5_W0_clk),
      // .W0_data(Mem5_W0_data)

      //W
      .clk0(Mem5_W0_clk),
      .csb0(~Mem5_W0_en),
      .addr0(Mem5_W0_addr),
      .din0(Mem5_W0_data),
      //R
      .clk1(Mem5_R0_clk),
      .csb1(1'b0),
      .addr1(Mem5_R0_addr),
      .dout1(Mem5_R0_data)
    );
    sram_128_256_scn4m_subm Mem6 ( // @[BuildingBlockNew.scala 39:25]
      // .R0_addr(Mem6_R0_addr),
      // .R0_clk(Mem6_R0_clk),
      // .R0_data(Mem6_R0_data),
      // .W0_addr(Mem6_W0_addr),
      // .W0_en(Mem6_W0_en),
      // .W0_clk(Mem6_W0_clk),
      // .W0_data(Mem6_W0_data)

      //W
      .clk0(Mem6_W0_clk),
      .csb0(~Mem6_W0_en),
      .addr0(Mem6_W0_addr),
      .din0(Mem6_W0_data),
      //R
      .clk1(Mem6_R0_clk),
      .csb1(1'b0),
      .addr1(Mem6_R0_addr),
      .dout1(Mem6_R0_data)
    );

  PEcol peCol ( // @[BuildingBlockNew.scala 83:21]
    .clock(peCol_clock),
    .reset(peCol_reset),
    .io_d_in_0_a(peCol_io_d_in_0_a),
    .io_d_in_0_valid_a(peCol_io_d_in_0_valid_a),
    .io_d_in_0_b(peCol_io_d_in_0_b),
    .io_d_in_1_a(peCol_io_d_in_1_a),
    .io_d_in_1_valid_a(peCol_io_d_in_1_valid_a),
    .io_d_in_1_b(peCol_io_d_in_1_b),
    .io_d_in_2_a(peCol_io_d_in_2_a),
    .io_d_in_2_valid_a(peCol_io_d_in_2_valid_a),
    .io_d_in_2_b(peCol_io_d_in_2_b),
    .io_d_in_3_a(peCol_io_d_in_3_a),
    .io_d_in_3_valid_a(peCol_io_d_in_3_valid_a),
    .io_d_in_3_b(peCol_io_d_in_3_b),
    .io_d_in_4_a(peCol_io_d_in_4_a),
    .io_d_in_4_valid_a(peCol_io_d_in_4_valid_a),
    .io_d_in_4_b(peCol_io_d_in_4_b),
    .io_d_in_5_a(peCol_io_d_in_5_a),
    .io_d_in_5_valid_a(peCol_io_d_in_5_valid_a),
    .io_d_in_5_b(peCol_io_d_in_5_b),
    .io_d_in_6_a(peCol_io_d_in_6_a),
    .io_d_in_6_valid_a(peCol_io_d_in_6_valid_a),
    .io_d_in_6_b(peCol_io_d_in_6_b),
    .io_d_in_7_a(peCol_io_d_in_7_a),
    .io_d_in_7_valid_a(peCol_io_d_in_7_valid_a),
    .io_d_in_7_b(peCol_io_d_in_7_b),
    .io_d_in_8_a(peCol_io_d_in_8_a),
    .io_d_in_8_valid_a(peCol_io_d_in_8_valid_a),
    .io_d_in_8_b(peCol_io_d_in_8_b),
    .io_d_in_9_a(peCol_io_d_in_9_a),
    .io_d_in_9_valid_a(peCol_io_d_in_9_valid_a),
    .io_d_in_9_b(peCol_io_d_in_9_b),
    .io_d_in_10_a(peCol_io_d_in_10_a),
    .io_d_in_10_valid_a(peCol_io_d_in_10_valid_a),
    .io_d_in_10_b(peCol_io_d_in_10_b),
    .io_d_in_11_a(peCol_io_d_in_11_a),
    .io_d_in_11_valid_a(peCol_io_d_in_11_valid_a),
    .io_d_in_11_b(peCol_io_d_in_11_b),
    .io_d_in_12_a(peCol_io_d_in_12_a),
    .io_d_in_12_valid_a(peCol_io_d_in_12_valid_a),
    .io_d_in_12_b(peCol_io_d_in_12_b),
    .io_d_in_13_a(peCol_io_d_in_13_a),
    .io_d_in_13_valid_a(peCol_io_d_in_13_valid_a),
    .io_d_in_13_b(peCol_io_d_in_13_b),
    .io_d_in_14_a(peCol_io_d_in_14_a),
    .io_d_in_14_valid_a(peCol_io_d_in_14_valid_a),
    .io_d_in_14_b(peCol_io_d_in_14_b),
    .io_d_in_15_a(peCol_io_d_in_15_a),
    .io_d_in_15_valid_a(peCol_io_d_in_15_valid_a),
    .io_d_in_15_b(peCol_io_d_in_15_b),
    .io_d_in_16_a(peCol_io_d_in_16_a),
    .io_d_in_16_valid_a(peCol_io_d_in_16_valid_a),
    .io_d_in_16_b(peCol_io_d_in_16_b),
    .io_d_in_17_a(peCol_io_d_in_17_a),
    .io_d_in_17_valid_a(peCol_io_d_in_17_valid_a),
    .io_d_in_17_b(peCol_io_d_in_17_b),
    .io_d_in_18_a(peCol_io_d_in_18_a),
    .io_d_in_18_valid_a(peCol_io_d_in_18_valid_a),
    .io_d_in_18_b(peCol_io_d_in_18_b),
    .io_d_in_19_a(peCol_io_d_in_19_a),
    .io_d_in_19_valid_a(peCol_io_d_in_19_valid_a),
    .io_d_in_19_b(peCol_io_d_in_19_b),
    .io_d_in_20_a(peCol_io_d_in_20_a),
    .io_d_in_20_valid_a(peCol_io_d_in_20_valid_a),
    .io_d_in_20_b(peCol_io_d_in_20_b),
    .io_d_in_21_a(peCol_io_d_in_21_a),
    .io_d_in_21_valid_a(peCol_io_d_in_21_valid_a),
    .io_d_in_21_b(peCol_io_d_in_21_b),
    .io_d_in_22_a(peCol_io_d_in_22_a),
    .io_d_in_22_valid_a(peCol_io_d_in_22_valid_a),
    .io_d_in_22_b(peCol_io_d_in_22_b),
    .io_d_in_23_a(peCol_io_d_in_23_a),
    .io_d_in_23_valid_a(peCol_io_d_in_23_valid_a),
    .io_d_in_23_b(peCol_io_d_in_23_b),
    .io_d_in_24_a(peCol_io_d_in_24_a),
    .io_d_in_24_valid_a(peCol_io_d_in_24_valid_a),
    .io_d_in_24_b(peCol_io_d_in_24_b),
    .io_d_in_25_a(peCol_io_d_in_25_a),
    .io_d_in_25_valid_a(peCol_io_d_in_25_valid_a),
    .io_d_in_25_b(peCol_io_d_in_25_b),
    .io_d_in_26_a(peCol_io_d_in_26_a),
    .io_d_in_26_valid_a(peCol_io_d_in_26_valid_a),
    .io_d_in_26_b(peCol_io_d_in_26_b),
    .io_d_in_27_a(peCol_io_d_in_27_a),
    .io_d_in_27_valid_a(peCol_io_d_in_27_valid_a),
    .io_d_in_27_b(peCol_io_d_in_27_b),
    .io_d_in_28_a(peCol_io_d_in_28_a),
    .io_d_in_28_valid_a(peCol_io_d_in_28_valid_a),
    .io_d_in_28_b(peCol_io_d_in_28_b),
    .io_d_in_29_a(peCol_io_d_in_29_a),
    .io_d_in_29_valid_a(peCol_io_d_in_29_valid_a),
    .io_d_in_29_b(peCol_io_d_in_29_b),
    .io_d_in_30_a(peCol_io_d_in_30_a),
    .io_d_in_30_valid_a(peCol_io_d_in_30_valid_a),
    .io_d_in_30_b(peCol_io_d_in_30_b),
    .io_d_in_31_a(peCol_io_d_in_31_a),
    .io_d_in_31_valid_a(peCol_io_d_in_31_valid_a),
    .io_d_in_31_b(peCol_io_d_in_31_b),
    .io_d_out_0_a(peCol_io_d_out_0_a),
    .io_d_out_0_valid_a(peCol_io_d_out_0_valid_a),
    .io_d_out_0_b(peCol_io_d_out_0_b),
    .io_d_out_1_a(peCol_io_d_out_1_a),
    .io_d_out_1_valid_a(peCol_io_d_out_1_valid_a),
    .io_d_out_1_b(peCol_io_d_out_1_b),
    .io_d_out_2_a(peCol_io_d_out_2_a),
    .io_d_out_2_valid_a(peCol_io_d_out_2_valid_a),
    .io_d_out_2_b(peCol_io_d_out_2_b),
    .io_d_out_3_a(peCol_io_d_out_3_a),
    .io_d_out_3_valid_a(peCol_io_d_out_3_valid_a),
    .io_d_out_3_b(peCol_io_d_out_3_b),
    .io_d_out_4_a(peCol_io_d_out_4_a),
    .io_d_out_4_valid_a(peCol_io_d_out_4_valid_a),
    .io_d_out_4_b(peCol_io_d_out_4_b),
    .io_d_out_5_a(peCol_io_d_out_5_a),
    .io_d_out_5_valid_a(peCol_io_d_out_5_valid_a),
    .io_d_out_5_b(peCol_io_d_out_5_b),
    .io_d_out_6_a(peCol_io_d_out_6_a),
    .io_d_out_6_valid_a(peCol_io_d_out_6_valid_a),
    .io_d_out_6_b(peCol_io_d_out_6_b),
    .io_d_out_7_a(peCol_io_d_out_7_a),
    .io_d_out_7_valid_a(peCol_io_d_out_7_valid_a),
    .io_d_out_7_b(peCol_io_d_out_7_b),
    .io_d_out_8_a(peCol_io_d_out_8_a),
    .io_d_out_8_valid_a(peCol_io_d_out_8_valid_a),
    .io_d_out_8_b(peCol_io_d_out_8_b),
    .io_d_out_9_a(peCol_io_d_out_9_a),
    .io_d_out_9_valid_a(peCol_io_d_out_9_valid_a),
    .io_d_out_9_b(peCol_io_d_out_9_b),
    .io_d_out_10_a(peCol_io_d_out_10_a),
    .io_d_out_10_valid_a(peCol_io_d_out_10_valid_a),
    .io_d_out_10_b(peCol_io_d_out_10_b),
    .io_d_out_11_a(peCol_io_d_out_11_a),
    .io_d_out_11_valid_a(peCol_io_d_out_11_valid_a),
    .io_d_out_11_b(peCol_io_d_out_11_b),
    .io_d_out_12_a(peCol_io_d_out_12_a),
    .io_d_out_12_valid_a(peCol_io_d_out_12_valid_a),
    .io_d_out_12_b(peCol_io_d_out_12_b),
    .io_d_out_13_a(peCol_io_d_out_13_a),
    .io_d_out_13_valid_a(peCol_io_d_out_13_valid_a),
    .io_d_out_13_b(peCol_io_d_out_13_b),
    .io_d_out_14_a(peCol_io_d_out_14_a),
    .io_d_out_14_valid_a(peCol_io_d_out_14_valid_a),
    .io_d_out_14_b(peCol_io_d_out_14_b),
    .io_d_out_15_a(peCol_io_d_out_15_a),
    .io_d_out_15_valid_a(peCol_io_d_out_15_valid_a),
    .io_d_out_15_b(peCol_io_d_out_15_b),
    .io_d_out_16_a(peCol_io_d_out_16_a),
    .io_d_out_16_valid_a(peCol_io_d_out_16_valid_a),
    .io_d_out_16_b(peCol_io_d_out_16_b),
    .io_d_out_17_a(peCol_io_d_out_17_a),
    .io_d_out_17_valid_a(peCol_io_d_out_17_valid_a),
    .io_d_out_17_b(peCol_io_d_out_17_b),
    .io_d_out_18_a(peCol_io_d_out_18_a),
    .io_d_out_18_valid_a(peCol_io_d_out_18_valid_a),
    .io_d_out_18_b(peCol_io_d_out_18_b),
    .io_d_out_19_a(peCol_io_d_out_19_a),
    .io_d_out_19_valid_a(peCol_io_d_out_19_valid_a),
    .io_d_out_19_b(peCol_io_d_out_19_b),
    .io_d_out_20_a(peCol_io_d_out_20_a),
    .io_d_out_20_valid_a(peCol_io_d_out_20_valid_a),
    .io_d_out_20_b(peCol_io_d_out_20_b),
    .io_d_out_21_a(peCol_io_d_out_21_a),
    .io_d_out_21_valid_a(peCol_io_d_out_21_valid_a),
    .io_d_out_21_b(peCol_io_d_out_21_b),
    .io_d_out_22_a(peCol_io_d_out_22_a),
    .io_d_out_22_valid_a(peCol_io_d_out_22_valid_a),
    .io_d_out_22_b(peCol_io_d_out_22_b),
    .io_d_out_23_a(peCol_io_d_out_23_a),
    .io_d_out_23_valid_a(peCol_io_d_out_23_valid_a),
    .io_d_out_23_b(peCol_io_d_out_23_b),
    .io_d_out_24_a(peCol_io_d_out_24_a),
    .io_d_out_24_valid_a(peCol_io_d_out_24_valid_a),
    .io_d_out_24_b(peCol_io_d_out_24_b),
    .io_d_out_25_a(peCol_io_d_out_25_a),
    .io_d_out_25_valid_a(peCol_io_d_out_25_valid_a),
    .io_d_out_25_b(peCol_io_d_out_25_b),
    .io_d_out_26_a(peCol_io_d_out_26_a),
    .io_d_out_26_valid_a(peCol_io_d_out_26_valid_a),
    .io_d_out_26_b(peCol_io_d_out_26_b),
    .io_d_out_27_a(peCol_io_d_out_27_a),
    .io_d_out_27_valid_a(peCol_io_d_out_27_valid_a),
    .io_d_out_27_b(peCol_io_d_out_27_b),
    .io_d_out_28_a(peCol_io_d_out_28_a),
    .io_d_out_28_valid_a(peCol_io_d_out_28_valid_a),
    .io_d_out_28_b(peCol_io_d_out_28_b),
    .io_d_out_29_a(peCol_io_d_out_29_a),
    .io_d_out_29_valid_a(peCol_io_d_out_29_valid_a),
    .io_d_out_29_b(peCol_io_d_out_29_b),
    .io_d_out_30_a(peCol_io_d_out_30_a),
    .io_d_out_30_valid_a(peCol_io_d_out_30_valid_a),
    .io_d_out_30_b(peCol_io_d_out_30_b),
    .io_d_out_31_a(peCol_io_d_out_31_a),
    .io_d_out_31_valid_a(peCol_io_d_out_31_valid_a),
    .io_d_out_31_b(peCol_io_d_out_31_b),
    .io_tagin_Tag(peCol_io_tagin_Tag),
    .io_tagin_RoundCnt(peCol_io_tagin_RoundCnt),
    .io_addrin(peCol_io_addrin),
    .io_tagout_Tag(peCol_io_tagout_Tag),
    .io_tagout_RoundCnt(peCol_io_tagout_RoundCnt),
    .io_addrout(peCol_io_addrout),
    .io_instr(peCol_io_instr)
  );
  CLOSingress1 ingress1 ( // @[BuildingBlockNew.scala 84:24]
    .clock(ingress1_clock),
    .io_in64_0(ingress1_io_in64_0),
    .io_in64_1(ingress1_io_in64_1),
    .io_in64_2(ingress1_io_in64_2),
    .io_in64_3(ingress1_io_in64_3),
    .io_in64_4(ingress1_io_in64_4),
    .io_in64_5(ingress1_io_in64_5),
    .io_in64_6(ingress1_io_in64_6),
    .io_in64_7(ingress1_io_in64_7),
    .io_in64_8(ingress1_io_in64_8),
    .io_in64_9(ingress1_io_in64_9),
    .io_in64_10(ingress1_io_in64_10),
    .io_in64_11(ingress1_io_in64_11),
    .io_in64_12(ingress1_io_in64_12),
    .io_in64_13(ingress1_io_in64_13),
    .io_in64_14(ingress1_io_in64_14),
    .io_in64_15(ingress1_io_in64_15),
    .io_in64_16(ingress1_io_in64_16),
    .io_in64_17(ingress1_io_in64_17),
    .io_in64_18(ingress1_io_in64_18),
    .io_in64_19(ingress1_io_in64_19),
    .io_in64_20(ingress1_io_in64_20),
    .io_in64_21(ingress1_io_in64_21),
    .io_in64_22(ingress1_io_in64_22),
    .io_in64_23(ingress1_io_in64_23),
    .io_in64_24(ingress1_io_in64_24),
    .io_in64_25(ingress1_io_in64_25),
    .io_in64_26(ingress1_io_in64_26),
    .io_in64_27(ingress1_io_in64_27),
    .io_in64_28(ingress1_io_in64_28),
    .io_in64_29(ingress1_io_in64_29),
    .io_in64_30(ingress1_io_in64_30),
    .io_in64_31(ingress1_io_in64_31),
    .io_in64_32(ingress1_io_in64_32),
    .io_in64_33(ingress1_io_in64_33),
    .io_in64_34(ingress1_io_in64_34),
    .io_in64_35(ingress1_io_in64_35),
    .io_in64_36(ingress1_io_in64_36),
    .io_in64_37(ingress1_io_in64_37),
    .io_in64_38(ingress1_io_in64_38),
    .io_in64_39(ingress1_io_in64_39),
    .io_in64_40(ingress1_io_in64_40),
    .io_in64_41(ingress1_io_in64_41),
    .io_in64_42(ingress1_io_in64_42),
    .io_in64_43(ingress1_io_in64_43),
    .io_in64_44(ingress1_io_in64_44),
    .io_in64_45(ingress1_io_in64_45),
    .io_in64_46(ingress1_io_in64_46),
    .io_in64_47(ingress1_io_in64_47),
    .io_in64_48(ingress1_io_in64_48),
    .io_in64_49(ingress1_io_in64_49),
    .io_in64_50(ingress1_io_in64_50),
    .io_in64_51(ingress1_io_in64_51),
    .io_in64_52(ingress1_io_in64_52),
    .io_in64_53(ingress1_io_in64_53),
    .io_in64_54(ingress1_io_in64_54),
    .io_in64_55(ingress1_io_in64_55),
    .io_in64_56(ingress1_io_in64_56),
    .io_in64_57(ingress1_io_in64_57),
    .io_in64_58(ingress1_io_in64_58),
    .io_in64_59(ingress1_io_in64_59),
    .io_in64_60(ingress1_io_in64_60),
    .io_in64_61(ingress1_io_in64_61),
    .io_in64_62(ingress1_io_in64_62),
    .io_in64_63(ingress1_io_in64_63),
    .io_validin64_0(ingress1_io_validin64_0),
    .io_validin64_2(ingress1_io_validin64_2),
    .io_validin64_4(ingress1_io_validin64_4),
    .io_validin64_6(ingress1_io_validin64_6),
    .io_validin64_8(ingress1_io_validin64_8),
    .io_validin64_10(ingress1_io_validin64_10),
    .io_validin64_12(ingress1_io_validin64_12),
    .io_validin64_14(ingress1_io_validin64_14),
    .io_validin64_16(ingress1_io_validin64_16),
    .io_validin64_18(ingress1_io_validin64_18),
    .io_validin64_20(ingress1_io_validin64_20),
    .io_validin64_22(ingress1_io_validin64_22),
    .io_validin64_24(ingress1_io_validin64_24),
    .io_validin64_26(ingress1_io_validin64_26),
    .io_validin64_28(ingress1_io_validin64_28),
    .io_validin64_30(ingress1_io_validin64_30),
    .io_validin64_32(ingress1_io_validin64_32),
    .io_validin64_34(ingress1_io_validin64_34),
    .io_validin64_36(ingress1_io_validin64_36),
    .io_validin64_38(ingress1_io_validin64_38),
    .io_validin64_40(ingress1_io_validin64_40),
    .io_validin64_42(ingress1_io_validin64_42),
    .io_validin64_44(ingress1_io_validin64_44),
    .io_validin64_46(ingress1_io_validin64_46),
    .io_validin64_48(ingress1_io_validin64_48),
    .io_validin64_50(ingress1_io_validin64_50),
    .io_validin64_52(ingress1_io_validin64_52),
    .io_validin64_54(ingress1_io_validin64_54),
    .io_validin64_56(ingress1_io_validin64_56),
    .io_validin64_58(ingress1_io_validin64_58),
    .io_validin64_60(ingress1_io_validin64_60),
    .io_validin64_62(ingress1_io_validin64_62),
    .io_tagin_Tag(ingress1_io_tagin_Tag),
    .io_tagin_RoundCnt(ingress1_io_tagin_RoundCnt),
    .io_addrin(ingress1_io_addrin),
    .io_out64_0(ingress1_io_out64_0),
    .io_out64_1(ingress1_io_out64_1),
    .io_out64_2(ingress1_io_out64_2),
    .io_out64_3(ingress1_io_out64_3),
    .io_out64_4(ingress1_io_out64_4),
    .io_out64_5(ingress1_io_out64_5),
    .io_out64_6(ingress1_io_out64_6),
    .io_out64_7(ingress1_io_out64_7),
    .io_out64_8(ingress1_io_out64_8),
    .io_out64_9(ingress1_io_out64_9),
    .io_out64_10(ingress1_io_out64_10),
    .io_out64_11(ingress1_io_out64_11),
    .io_out64_12(ingress1_io_out64_12),
    .io_out64_13(ingress1_io_out64_13),
    .io_out64_14(ingress1_io_out64_14),
    .io_out64_15(ingress1_io_out64_15),
    .io_out64_16(ingress1_io_out64_16),
    .io_out64_17(ingress1_io_out64_17),
    .io_out64_18(ingress1_io_out64_18),
    .io_out64_19(ingress1_io_out64_19),
    .io_out64_20(ingress1_io_out64_20),
    .io_out64_21(ingress1_io_out64_21),
    .io_out64_22(ingress1_io_out64_22),
    .io_out64_23(ingress1_io_out64_23),
    .io_out64_24(ingress1_io_out64_24),
    .io_out64_25(ingress1_io_out64_25),
    .io_out64_26(ingress1_io_out64_26),
    .io_out64_27(ingress1_io_out64_27),
    .io_out64_28(ingress1_io_out64_28),
    .io_out64_29(ingress1_io_out64_29),
    .io_out64_30(ingress1_io_out64_30),
    .io_out64_31(ingress1_io_out64_31),
    .io_out64_32(ingress1_io_out64_32),
    .io_out64_33(ingress1_io_out64_33),
    .io_out64_34(ingress1_io_out64_34),
    .io_out64_35(ingress1_io_out64_35),
    .io_out64_36(ingress1_io_out64_36),
    .io_out64_37(ingress1_io_out64_37),
    .io_out64_38(ingress1_io_out64_38),
    .io_out64_39(ingress1_io_out64_39),
    .io_out64_40(ingress1_io_out64_40),
    .io_out64_41(ingress1_io_out64_41),
    .io_out64_42(ingress1_io_out64_42),
    .io_out64_43(ingress1_io_out64_43),
    .io_out64_44(ingress1_io_out64_44),
    .io_out64_45(ingress1_io_out64_45),
    .io_out64_46(ingress1_io_out64_46),
    .io_out64_47(ingress1_io_out64_47),
    .io_out64_48(ingress1_io_out64_48),
    .io_out64_49(ingress1_io_out64_49),
    .io_out64_50(ingress1_io_out64_50),
    .io_out64_51(ingress1_io_out64_51),
    .io_out64_52(ingress1_io_out64_52),
    .io_out64_53(ingress1_io_out64_53),
    .io_out64_54(ingress1_io_out64_54),
    .io_out64_55(ingress1_io_out64_55),
    .io_out64_56(ingress1_io_out64_56),
    .io_out64_57(ingress1_io_out64_57),
    .io_out64_58(ingress1_io_out64_58),
    .io_out64_59(ingress1_io_out64_59),
    .io_out64_60(ingress1_io_out64_60),
    .io_out64_61(ingress1_io_out64_61),
    .io_out64_62(ingress1_io_out64_62),
    .io_out64_63(ingress1_io_out64_63),
    .io_validout64_0(ingress1_io_validout64_0),
    .io_validout64_1(ingress1_io_validout64_1),
    .io_validout64_2(ingress1_io_validout64_2),
    .io_validout64_3(ingress1_io_validout64_3),
    .io_validout64_4(ingress1_io_validout64_4),
    .io_validout64_5(ingress1_io_validout64_5),
    .io_validout64_6(ingress1_io_validout64_6),
    .io_validout64_7(ingress1_io_validout64_7),
    .io_validout64_8(ingress1_io_validout64_8),
    .io_validout64_9(ingress1_io_validout64_9),
    .io_validout64_10(ingress1_io_validout64_10),
    .io_validout64_11(ingress1_io_validout64_11),
    .io_validout64_12(ingress1_io_validout64_12),
    .io_validout64_13(ingress1_io_validout64_13),
    .io_validout64_14(ingress1_io_validout64_14),
    .io_validout64_15(ingress1_io_validout64_15),
    .io_validout64_16(ingress1_io_validout64_16),
    .io_validout64_17(ingress1_io_validout64_17),
    .io_validout64_18(ingress1_io_validout64_18),
    .io_validout64_19(ingress1_io_validout64_19),
    .io_validout64_20(ingress1_io_validout64_20),
    .io_validout64_21(ingress1_io_validout64_21),
    .io_validout64_22(ingress1_io_validout64_22),
    .io_validout64_23(ingress1_io_validout64_23),
    .io_validout64_24(ingress1_io_validout64_24),
    .io_validout64_25(ingress1_io_validout64_25),
    .io_validout64_26(ingress1_io_validout64_26),
    .io_validout64_27(ingress1_io_validout64_27),
    .io_validout64_28(ingress1_io_validout64_28),
    .io_validout64_29(ingress1_io_validout64_29),
    .io_validout64_30(ingress1_io_validout64_30),
    .io_validout64_31(ingress1_io_validout64_31),
    .io_validout64_32(ingress1_io_validout64_32),
    .io_validout64_33(ingress1_io_validout64_33),
    .io_validout64_34(ingress1_io_validout64_34),
    .io_validout64_35(ingress1_io_validout64_35),
    .io_validout64_36(ingress1_io_validout64_36),
    .io_validout64_37(ingress1_io_validout64_37),
    .io_validout64_38(ingress1_io_validout64_38),
    .io_validout64_39(ingress1_io_validout64_39),
    .io_validout64_40(ingress1_io_validout64_40),
    .io_validout64_41(ingress1_io_validout64_41),
    .io_validout64_42(ingress1_io_validout64_42),
    .io_validout64_43(ingress1_io_validout64_43),
    .io_validout64_44(ingress1_io_validout64_44),
    .io_validout64_45(ingress1_io_validout64_45),
    .io_validout64_46(ingress1_io_validout64_46),
    .io_validout64_47(ingress1_io_validout64_47),
    .io_validout64_48(ingress1_io_validout64_48),
    .io_validout64_49(ingress1_io_validout64_49),
    .io_validout64_50(ingress1_io_validout64_50),
    .io_validout64_51(ingress1_io_validout64_51),
    .io_validout64_52(ingress1_io_validout64_52),
    .io_validout64_53(ingress1_io_validout64_53),
    .io_validout64_54(ingress1_io_validout64_54),
    .io_validout64_55(ingress1_io_validout64_55),
    .io_validout64_56(ingress1_io_validout64_56),
    .io_validout64_57(ingress1_io_validout64_57),
    .io_validout64_58(ingress1_io_validout64_58),
    .io_validout64_59(ingress1_io_validout64_59),
    .io_validout64_60(ingress1_io_validout64_60),
    .io_validout64_61(ingress1_io_validout64_61),
    .io_validout64_62(ingress1_io_validout64_62),
    .io_validout64_63(ingress1_io_validout64_63),
    .io_tagout_Tag(ingress1_io_tagout_Tag),
    .io_tagout_RoundCnt(ingress1_io_tagout_RoundCnt),
    .io_addrout(ingress1_io_addrout),
    .io_ctrl(ingress1_io_ctrl)
  );
  CLOSingress2 ingress2 ( // @[BuildingBlockNew.scala 85:24]
    .clock(ingress2_clock),
    .io_in64_0(ingress2_io_in64_0),
    .io_in64_1(ingress2_io_in64_1),
    .io_in64_2(ingress2_io_in64_2),
    .io_in64_3(ingress2_io_in64_3),
    .io_in64_4(ingress2_io_in64_4),
    .io_in64_5(ingress2_io_in64_5),
    .io_in64_6(ingress2_io_in64_6),
    .io_in64_7(ingress2_io_in64_7),
    .io_in64_8(ingress2_io_in64_8),
    .io_in64_9(ingress2_io_in64_9),
    .io_in64_10(ingress2_io_in64_10),
    .io_in64_11(ingress2_io_in64_11),
    .io_in64_12(ingress2_io_in64_12),
    .io_in64_13(ingress2_io_in64_13),
    .io_in64_14(ingress2_io_in64_14),
    .io_in64_15(ingress2_io_in64_15),
    .io_in64_16(ingress2_io_in64_16),
    .io_in64_17(ingress2_io_in64_17),
    .io_in64_18(ingress2_io_in64_18),
    .io_in64_19(ingress2_io_in64_19),
    .io_in64_20(ingress2_io_in64_20),
    .io_in64_21(ingress2_io_in64_21),
    .io_in64_22(ingress2_io_in64_22),
    .io_in64_23(ingress2_io_in64_23),
    .io_in64_24(ingress2_io_in64_24),
    .io_in64_25(ingress2_io_in64_25),
    .io_in64_26(ingress2_io_in64_26),
    .io_in64_27(ingress2_io_in64_27),
    .io_in64_28(ingress2_io_in64_28),
    .io_in64_29(ingress2_io_in64_29),
    .io_in64_30(ingress2_io_in64_30),
    .io_in64_31(ingress2_io_in64_31),
    .io_in64_32(ingress2_io_in64_32),
    .io_in64_33(ingress2_io_in64_33),
    .io_in64_34(ingress2_io_in64_34),
    .io_in64_35(ingress2_io_in64_35),
    .io_in64_36(ingress2_io_in64_36),
    .io_in64_37(ingress2_io_in64_37),
    .io_in64_38(ingress2_io_in64_38),
    .io_in64_39(ingress2_io_in64_39),
    .io_in64_40(ingress2_io_in64_40),
    .io_in64_41(ingress2_io_in64_41),
    .io_in64_42(ingress2_io_in64_42),
    .io_in64_43(ingress2_io_in64_43),
    .io_in64_44(ingress2_io_in64_44),
    .io_in64_45(ingress2_io_in64_45),
    .io_in64_46(ingress2_io_in64_46),
    .io_in64_47(ingress2_io_in64_47),
    .io_in64_48(ingress2_io_in64_48),
    .io_in64_49(ingress2_io_in64_49),
    .io_in64_50(ingress2_io_in64_50),
    .io_in64_51(ingress2_io_in64_51),
    .io_in64_52(ingress2_io_in64_52),
    .io_in64_53(ingress2_io_in64_53),
    .io_in64_54(ingress2_io_in64_54),
    .io_in64_55(ingress2_io_in64_55),
    .io_in64_56(ingress2_io_in64_56),
    .io_in64_57(ingress2_io_in64_57),
    .io_in64_58(ingress2_io_in64_58),
    .io_in64_59(ingress2_io_in64_59),
    .io_in64_60(ingress2_io_in64_60),
    .io_in64_61(ingress2_io_in64_61),
    .io_in64_62(ingress2_io_in64_62),
    .io_in64_63(ingress2_io_in64_63),
    .io_validin64_0(ingress2_io_validin64_0),
    .io_validin64_1(ingress2_io_validin64_1),
    .io_validin64_2(ingress2_io_validin64_2),
    .io_validin64_3(ingress2_io_validin64_3),
    .io_validin64_4(ingress2_io_validin64_4),
    .io_validin64_5(ingress2_io_validin64_5),
    .io_validin64_6(ingress2_io_validin64_6),
    .io_validin64_7(ingress2_io_validin64_7),
    .io_validin64_8(ingress2_io_validin64_8),
    .io_validin64_9(ingress2_io_validin64_9),
    .io_validin64_10(ingress2_io_validin64_10),
    .io_validin64_11(ingress2_io_validin64_11),
    .io_validin64_12(ingress2_io_validin64_12),
    .io_validin64_13(ingress2_io_validin64_13),
    .io_validin64_14(ingress2_io_validin64_14),
    .io_validin64_15(ingress2_io_validin64_15),
    .io_validin64_16(ingress2_io_validin64_16),
    .io_validin64_17(ingress2_io_validin64_17),
    .io_validin64_18(ingress2_io_validin64_18),
    .io_validin64_19(ingress2_io_validin64_19),
    .io_validin64_20(ingress2_io_validin64_20),
    .io_validin64_21(ingress2_io_validin64_21),
    .io_validin64_22(ingress2_io_validin64_22),
    .io_validin64_23(ingress2_io_validin64_23),
    .io_validin64_24(ingress2_io_validin64_24),
    .io_validin64_25(ingress2_io_validin64_25),
    .io_validin64_26(ingress2_io_validin64_26),
    .io_validin64_27(ingress2_io_validin64_27),
    .io_validin64_28(ingress2_io_validin64_28),
    .io_validin64_29(ingress2_io_validin64_29),
    .io_validin64_30(ingress2_io_validin64_30),
    .io_validin64_31(ingress2_io_validin64_31),
    .io_validin64_32(ingress2_io_validin64_32),
    .io_validin64_33(ingress2_io_validin64_33),
    .io_validin64_34(ingress2_io_validin64_34),
    .io_validin64_35(ingress2_io_validin64_35),
    .io_validin64_36(ingress2_io_validin64_36),
    .io_validin64_37(ingress2_io_validin64_37),
    .io_validin64_38(ingress2_io_validin64_38),
    .io_validin64_39(ingress2_io_validin64_39),
    .io_validin64_40(ingress2_io_validin64_40),
    .io_validin64_41(ingress2_io_validin64_41),
    .io_validin64_42(ingress2_io_validin64_42),
    .io_validin64_43(ingress2_io_validin64_43),
    .io_validin64_44(ingress2_io_validin64_44),
    .io_validin64_45(ingress2_io_validin64_45),
    .io_validin64_46(ingress2_io_validin64_46),
    .io_validin64_47(ingress2_io_validin64_47),
    .io_validin64_48(ingress2_io_validin64_48),
    .io_validin64_49(ingress2_io_validin64_49),
    .io_validin64_50(ingress2_io_validin64_50),
    .io_validin64_51(ingress2_io_validin64_51),
    .io_validin64_52(ingress2_io_validin64_52),
    .io_validin64_53(ingress2_io_validin64_53),
    .io_validin64_54(ingress2_io_validin64_54),
    .io_validin64_55(ingress2_io_validin64_55),
    .io_validin64_56(ingress2_io_validin64_56),
    .io_validin64_57(ingress2_io_validin64_57),
    .io_validin64_58(ingress2_io_validin64_58),
    .io_validin64_59(ingress2_io_validin64_59),
    .io_validin64_60(ingress2_io_validin64_60),
    .io_validin64_61(ingress2_io_validin64_61),
    .io_validin64_62(ingress2_io_validin64_62),
    .io_validin64_63(ingress2_io_validin64_63),
    .io_tagin_Tag(ingress2_io_tagin_Tag),
    .io_tagin_RoundCnt(ingress2_io_tagin_RoundCnt),
    .io_addrin(ingress2_io_addrin),
    .io_out64_0(ingress2_io_out64_0),
    .io_out64_1(ingress2_io_out64_1),
    .io_out64_2(ingress2_io_out64_2),
    .io_out64_3(ingress2_io_out64_3),
    .io_out64_4(ingress2_io_out64_4),
    .io_out64_5(ingress2_io_out64_5),
    .io_out64_6(ingress2_io_out64_6),
    .io_out64_7(ingress2_io_out64_7),
    .io_out64_8(ingress2_io_out64_8),
    .io_out64_9(ingress2_io_out64_9),
    .io_out64_10(ingress2_io_out64_10),
    .io_out64_11(ingress2_io_out64_11),
    .io_out64_12(ingress2_io_out64_12),
    .io_out64_13(ingress2_io_out64_13),
    .io_out64_14(ingress2_io_out64_14),
    .io_out64_15(ingress2_io_out64_15),
    .io_out64_16(ingress2_io_out64_16),
    .io_out64_17(ingress2_io_out64_17),
    .io_out64_18(ingress2_io_out64_18),
    .io_out64_19(ingress2_io_out64_19),
    .io_out64_20(ingress2_io_out64_20),
    .io_out64_21(ingress2_io_out64_21),
    .io_out64_22(ingress2_io_out64_22),
    .io_out64_23(ingress2_io_out64_23),
    .io_out64_24(ingress2_io_out64_24),
    .io_out64_25(ingress2_io_out64_25),
    .io_out64_26(ingress2_io_out64_26),
    .io_out64_27(ingress2_io_out64_27),
    .io_out64_28(ingress2_io_out64_28),
    .io_out64_29(ingress2_io_out64_29),
    .io_out64_30(ingress2_io_out64_30),
    .io_out64_31(ingress2_io_out64_31),
    .io_out64_32(ingress2_io_out64_32),
    .io_out64_33(ingress2_io_out64_33),
    .io_out64_34(ingress2_io_out64_34),
    .io_out64_35(ingress2_io_out64_35),
    .io_out64_36(ingress2_io_out64_36),
    .io_out64_37(ingress2_io_out64_37),
    .io_out64_38(ingress2_io_out64_38),
    .io_out64_39(ingress2_io_out64_39),
    .io_out64_40(ingress2_io_out64_40),
    .io_out64_41(ingress2_io_out64_41),
    .io_out64_42(ingress2_io_out64_42),
    .io_out64_43(ingress2_io_out64_43),
    .io_out64_44(ingress2_io_out64_44),
    .io_out64_45(ingress2_io_out64_45),
    .io_out64_46(ingress2_io_out64_46),
    .io_out64_47(ingress2_io_out64_47),
    .io_out64_48(ingress2_io_out64_48),
    .io_out64_49(ingress2_io_out64_49),
    .io_out64_50(ingress2_io_out64_50),
    .io_out64_51(ingress2_io_out64_51),
    .io_out64_52(ingress2_io_out64_52),
    .io_out64_53(ingress2_io_out64_53),
    .io_out64_54(ingress2_io_out64_54),
    .io_out64_55(ingress2_io_out64_55),
    .io_out64_56(ingress2_io_out64_56),
    .io_out64_57(ingress2_io_out64_57),
    .io_out64_58(ingress2_io_out64_58),
    .io_out64_59(ingress2_io_out64_59),
    .io_out64_60(ingress2_io_out64_60),
    .io_out64_61(ingress2_io_out64_61),
    .io_out64_62(ingress2_io_out64_62),
    .io_out64_63(ingress2_io_out64_63),
    .io_validout64_0(ingress2_io_validout64_0),
    .io_validout64_1(ingress2_io_validout64_1),
    .io_validout64_2(ingress2_io_validout64_2),
    .io_validout64_3(ingress2_io_validout64_3),
    .io_validout64_4(ingress2_io_validout64_4),
    .io_validout64_5(ingress2_io_validout64_5),
    .io_validout64_6(ingress2_io_validout64_6),
    .io_validout64_7(ingress2_io_validout64_7),
    .io_validout64_8(ingress2_io_validout64_8),
    .io_validout64_9(ingress2_io_validout64_9),
    .io_validout64_10(ingress2_io_validout64_10),
    .io_validout64_11(ingress2_io_validout64_11),
    .io_validout64_12(ingress2_io_validout64_12),
    .io_validout64_13(ingress2_io_validout64_13),
    .io_validout64_14(ingress2_io_validout64_14),
    .io_validout64_15(ingress2_io_validout64_15),
    .io_validout64_16(ingress2_io_validout64_16),
    .io_validout64_17(ingress2_io_validout64_17),
    .io_validout64_18(ingress2_io_validout64_18),
    .io_validout64_19(ingress2_io_validout64_19),
    .io_validout64_20(ingress2_io_validout64_20),
    .io_validout64_21(ingress2_io_validout64_21),
    .io_validout64_22(ingress2_io_validout64_22),
    .io_validout64_23(ingress2_io_validout64_23),
    .io_validout64_24(ingress2_io_validout64_24),
    .io_validout64_25(ingress2_io_validout64_25),
    .io_validout64_26(ingress2_io_validout64_26),
    .io_validout64_27(ingress2_io_validout64_27),
    .io_validout64_28(ingress2_io_validout64_28),
    .io_validout64_29(ingress2_io_validout64_29),
    .io_validout64_30(ingress2_io_validout64_30),
    .io_validout64_31(ingress2_io_validout64_31),
    .io_validout64_32(ingress2_io_validout64_32),
    .io_validout64_33(ingress2_io_validout64_33),
    .io_validout64_34(ingress2_io_validout64_34),
    .io_validout64_35(ingress2_io_validout64_35),
    .io_validout64_36(ingress2_io_validout64_36),
    .io_validout64_37(ingress2_io_validout64_37),
    .io_validout64_38(ingress2_io_validout64_38),
    .io_validout64_39(ingress2_io_validout64_39),
    .io_validout64_40(ingress2_io_validout64_40),
    .io_validout64_41(ingress2_io_validout64_41),
    .io_validout64_42(ingress2_io_validout64_42),
    .io_validout64_43(ingress2_io_validout64_43),
    .io_validout64_44(ingress2_io_validout64_44),
    .io_validout64_45(ingress2_io_validout64_45),
    .io_validout64_46(ingress2_io_validout64_46),
    .io_validout64_47(ingress2_io_validout64_47),
    .io_validout64_48(ingress2_io_validout64_48),
    .io_validout64_49(ingress2_io_validout64_49),
    .io_validout64_50(ingress2_io_validout64_50),
    .io_validout64_51(ingress2_io_validout64_51),
    .io_validout64_52(ingress2_io_validout64_52),
    .io_validout64_53(ingress2_io_validout64_53),
    .io_validout64_54(ingress2_io_validout64_54),
    .io_validout64_55(ingress2_io_validout64_55),
    .io_validout64_56(ingress2_io_validout64_56),
    .io_validout64_57(ingress2_io_validout64_57),
    .io_validout64_58(ingress2_io_validout64_58),
    .io_validout64_59(ingress2_io_validout64_59),
    .io_validout64_60(ingress2_io_validout64_60),
    .io_validout64_61(ingress2_io_validout64_61),
    .io_validout64_62(ingress2_io_validout64_62),
    .io_validout64_63(ingress2_io_validout64_63),
    .io_tagout_Tag(ingress2_io_tagout_Tag),
    .io_tagout_RoundCnt(ingress2_io_tagout_RoundCnt),
    .io_addrout(ingress2_io_addrout),
    .io_ctrl(ingress2_io_ctrl)
  );
  CLOSingress2 middle ( // @[BuildingBlockNew.scala 86:22]
    .clock(middle_clock),
    .io_in64_0(middle_io_in64_0),
    .io_in64_1(middle_io_in64_1),
    .io_in64_2(middle_io_in64_2),
    .io_in64_3(middle_io_in64_3),
    .io_in64_4(middle_io_in64_4),
    .io_in64_5(middle_io_in64_5),
    .io_in64_6(middle_io_in64_6),
    .io_in64_7(middle_io_in64_7),
    .io_in64_8(middle_io_in64_8),
    .io_in64_9(middle_io_in64_9),
    .io_in64_10(middle_io_in64_10),
    .io_in64_11(middle_io_in64_11),
    .io_in64_12(middle_io_in64_12),
    .io_in64_13(middle_io_in64_13),
    .io_in64_14(middle_io_in64_14),
    .io_in64_15(middle_io_in64_15),
    .io_in64_16(middle_io_in64_16),
    .io_in64_17(middle_io_in64_17),
    .io_in64_18(middle_io_in64_18),
    .io_in64_19(middle_io_in64_19),
    .io_in64_20(middle_io_in64_20),
    .io_in64_21(middle_io_in64_21),
    .io_in64_22(middle_io_in64_22),
    .io_in64_23(middle_io_in64_23),
    .io_in64_24(middle_io_in64_24),
    .io_in64_25(middle_io_in64_25),
    .io_in64_26(middle_io_in64_26),
    .io_in64_27(middle_io_in64_27),
    .io_in64_28(middle_io_in64_28),
    .io_in64_29(middle_io_in64_29),
    .io_in64_30(middle_io_in64_30),
    .io_in64_31(middle_io_in64_31),
    .io_in64_32(middle_io_in64_32),
    .io_in64_33(middle_io_in64_33),
    .io_in64_34(middle_io_in64_34),
    .io_in64_35(middle_io_in64_35),
    .io_in64_36(middle_io_in64_36),
    .io_in64_37(middle_io_in64_37),
    .io_in64_38(middle_io_in64_38),
    .io_in64_39(middle_io_in64_39),
    .io_in64_40(middle_io_in64_40),
    .io_in64_41(middle_io_in64_41),
    .io_in64_42(middle_io_in64_42),
    .io_in64_43(middle_io_in64_43),
    .io_in64_44(middle_io_in64_44),
    .io_in64_45(middle_io_in64_45),
    .io_in64_46(middle_io_in64_46),
    .io_in64_47(middle_io_in64_47),
    .io_in64_48(middle_io_in64_48),
    .io_in64_49(middle_io_in64_49),
    .io_in64_50(middle_io_in64_50),
    .io_in64_51(middle_io_in64_51),
    .io_in64_52(middle_io_in64_52),
    .io_in64_53(middle_io_in64_53),
    .io_in64_54(middle_io_in64_54),
    .io_in64_55(middle_io_in64_55),
    .io_in64_56(middle_io_in64_56),
    .io_in64_57(middle_io_in64_57),
    .io_in64_58(middle_io_in64_58),
    .io_in64_59(middle_io_in64_59),
    .io_in64_60(middle_io_in64_60),
    .io_in64_61(middle_io_in64_61),
    .io_in64_62(middle_io_in64_62),
    .io_in64_63(middle_io_in64_63),
    .io_validin64_0(middle_io_validin64_0),
    .io_validin64_1(middle_io_validin64_1),
    .io_validin64_2(middle_io_validin64_2),
    .io_validin64_3(middle_io_validin64_3),
    .io_validin64_4(middle_io_validin64_4),
    .io_validin64_5(middle_io_validin64_5),
    .io_validin64_6(middle_io_validin64_6),
    .io_validin64_7(middle_io_validin64_7),
    .io_validin64_8(middle_io_validin64_8),
    .io_validin64_9(middle_io_validin64_9),
    .io_validin64_10(middle_io_validin64_10),
    .io_validin64_11(middle_io_validin64_11),
    .io_validin64_12(middle_io_validin64_12),
    .io_validin64_13(middle_io_validin64_13),
    .io_validin64_14(middle_io_validin64_14),
    .io_validin64_15(middle_io_validin64_15),
    .io_validin64_16(middle_io_validin64_16),
    .io_validin64_17(middle_io_validin64_17),
    .io_validin64_18(middle_io_validin64_18),
    .io_validin64_19(middle_io_validin64_19),
    .io_validin64_20(middle_io_validin64_20),
    .io_validin64_21(middle_io_validin64_21),
    .io_validin64_22(middle_io_validin64_22),
    .io_validin64_23(middle_io_validin64_23),
    .io_validin64_24(middle_io_validin64_24),
    .io_validin64_25(middle_io_validin64_25),
    .io_validin64_26(middle_io_validin64_26),
    .io_validin64_27(middle_io_validin64_27),
    .io_validin64_28(middle_io_validin64_28),
    .io_validin64_29(middle_io_validin64_29),
    .io_validin64_30(middle_io_validin64_30),
    .io_validin64_31(middle_io_validin64_31),
    .io_validin64_32(middle_io_validin64_32),
    .io_validin64_33(middle_io_validin64_33),
    .io_validin64_34(middle_io_validin64_34),
    .io_validin64_35(middle_io_validin64_35),
    .io_validin64_36(middle_io_validin64_36),
    .io_validin64_37(middle_io_validin64_37),
    .io_validin64_38(middle_io_validin64_38),
    .io_validin64_39(middle_io_validin64_39),
    .io_validin64_40(middle_io_validin64_40),
    .io_validin64_41(middle_io_validin64_41),
    .io_validin64_42(middle_io_validin64_42),
    .io_validin64_43(middle_io_validin64_43),
    .io_validin64_44(middle_io_validin64_44),
    .io_validin64_45(middle_io_validin64_45),
    .io_validin64_46(middle_io_validin64_46),
    .io_validin64_47(middle_io_validin64_47),
    .io_validin64_48(middle_io_validin64_48),
    .io_validin64_49(middle_io_validin64_49),
    .io_validin64_50(middle_io_validin64_50),
    .io_validin64_51(middle_io_validin64_51),
    .io_validin64_52(middle_io_validin64_52),
    .io_validin64_53(middle_io_validin64_53),
    .io_validin64_54(middle_io_validin64_54),
    .io_validin64_55(middle_io_validin64_55),
    .io_validin64_56(middle_io_validin64_56),
    .io_validin64_57(middle_io_validin64_57),
    .io_validin64_58(middle_io_validin64_58),
    .io_validin64_59(middle_io_validin64_59),
    .io_validin64_60(middle_io_validin64_60),
    .io_validin64_61(middle_io_validin64_61),
    .io_validin64_62(middle_io_validin64_62),
    .io_validin64_63(middle_io_validin64_63),
    .io_tagin_Tag(middle_io_tagin_Tag),
    .io_tagin_RoundCnt(middle_io_tagin_RoundCnt),
    .io_addrin(middle_io_addrin),
    .io_out64_0(middle_io_out64_0),
    .io_out64_1(middle_io_out64_1),
    .io_out64_2(middle_io_out64_2),
    .io_out64_3(middle_io_out64_3),
    .io_out64_4(middle_io_out64_4),
    .io_out64_5(middle_io_out64_5),
    .io_out64_6(middle_io_out64_6),
    .io_out64_7(middle_io_out64_7),
    .io_out64_8(middle_io_out64_8),
    .io_out64_9(middle_io_out64_9),
    .io_out64_10(middle_io_out64_10),
    .io_out64_11(middle_io_out64_11),
    .io_out64_12(middle_io_out64_12),
    .io_out64_13(middle_io_out64_13),
    .io_out64_14(middle_io_out64_14),
    .io_out64_15(middle_io_out64_15),
    .io_out64_16(middle_io_out64_16),
    .io_out64_17(middle_io_out64_17),
    .io_out64_18(middle_io_out64_18),
    .io_out64_19(middle_io_out64_19),
    .io_out64_20(middle_io_out64_20),
    .io_out64_21(middle_io_out64_21),
    .io_out64_22(middle_io_out64_22),
    .io_out64_23(middle_io_out64_23),
    .io_out64_24(middle_io_out64_24),
    .io_out64_25(middle_io_out64_25),
    .io_out64_26(middle_io_out64_26),
    .io_out64_27(middle_io_out64_27),
    .io_out64_28(middle_io_out64_28),
    .io_out64_29(middle_io_out64_29),
    .io_out64_30(middle_io_out64_30),
    .io_out64_31(middle_io_out64_31),
    .io_out64_32(middle_io_out64_32),
    .io_out64_33(middle_io_out64_33),
    .io_out64_34(middle_io_out64_34),
    .io_out64_35(middle_io_out64_35),
    .io_out64_36(middle_io_out64_36),
    .io_out64_37(middle_io_out64_37),
    .io_out64_38(middle_io_out64_38),
    .io_out64_39(middle_io_out64_39),
    .io_out64_40(middle_io_out64_40),
    .io_out64_41(middle_io_out64_41),
    .io_out64_42(middle_io_out64_42),
    .io_out64_43(middle_io_out64_43),
    .io_out64_44(middle_io_out64_44),
    .io_out64_45(middle_io_out64_45),
    .io_out64_46(middle_io_out64_46),
    .io_out64_47(middle_io_out64_47),
    .io_out64_48(middle_io_out64_48),
    .io_out64_49(middle_io_out64_49),
    .io_out64_50(middle_io_out64_50),
    .io_out64_51(middle_io_out64_51),
    .io_out64_52(middle_io_out64_52),
    .io_out64_53(middle_io_out64_53),
    .io_out64_54(middle_io_out64_54),
    .io_out64_55(middle_io_out64_55),
    .io_out64_56(middle_io_out64_56),
    .io_out64_57(middle_io_out64_57),
    .io_out64_58(middle_io_out64_58),
    .io_out64_59(middle_io_out64_59),
    .io_out64_60(middle_io_out64_60),
    .io_out64_61(middle_io_out64_61),
    .io_out64_62(middle_io_out64_62),
    .io_out64_63(middle_io_out64_63),
    .io_validout64_0(middle_io_validout64_0),
    .io_validout64_1(middle_io_validout64_1),
    .io_validout64_2(middle_io_validout64_2),
    .io_validout64_3(middle_io_validout64_3),
    .io_validout64_4(middle_io_validout64_4),
    .io_validout64_5(middle_io_validout64_5),
    .io_validout64_6(middle_io_validout64_6),
    .io_validout64_7(middle_io_validout64_7),
    .io_validout64_8(middle_io_validout64_8),
    .io_validout64_9(middle_io_validout64_9),
    .io_validout64_10(middle_io_validout64_10),
    .io_validout64_11(middle_io_validout64_11),
    .io_validout64_12(middle_io_validout64_12),
    .io_validout64_13(middle_io_validout64_13),
    .io_validout64_14(middle_io_validout64_14),
    .io_validout64_15(middle_io_validout64_15),
    .io_validout64_16(middle_io_validout64_16),
    .io_validout64_17(middle_io_validout64_17),
    .io_validout64_18(middle_io_validout64_18),
    .io_validout64_19(middle_io_validout64_19),
    .io_validout64_20(middle_io_validout64_20),
    .io_validout64_21(middle_io_validout64_21),
    .io_validout64_22(middle_io_validout64_22),
    .io_validout64_23(middle_io_validout64_23),
    .io_validout64_24(middle_io_validout64_24),
    .io_validout64_25(middle_io_validout64_25),
    .io_validout64_26(middle_io_validout64_26),
    .io_validout64_27(middle_io_validout64_27),
    .io_validout64_28(middle_io_validout64_28),
    .io_validout64_29(middle_io_validout64_29),
    .io_validout64_30(middle_io_validout64_30),
    .io_validout64_31(middle_io_validout64_31),
    .io_validout64_32(middle_io_validout64_32),
    .io_validout64_33(middle_io_validout64_33),
    .io_validout64_34(middle_io_validout64_34),
    .io_validout64_35(middle_io_validout64_35),
    .io_validout64_36(middle_io_validout64_36),
    .io_validout64_37(middle_io_validout64_37),
    .io_validout64_38(middle_io_validout64_38),
    .io_validout64_39(middle_io_validout64_39),
    .io_validout64_40(middle_io_validout64_40),
    .io_validout64_41(middle_io_validout64_41),
    .io_validout64_42(middle_io_validout64_42),
    .io_validout64_43(middle_io_validout64_43),
    .io_validout64_44(middle_io_validout64_44),
    .io_validout64_45(middle_io_validout64_45),
    .io_validout64_46(middle_io_validout64_46),
    .io_validout64_47(middle_io_validout64_47),
    .io_validout64_48(middle_io_validout64_48),
    .io_validout64_49(middle_io_validout64_49),
    .io_validout64_50(middle_io_validout64_50),
    .io_validout64_51(middle_io_validout64_51),
    .io_validout64_52(middle_io_validout64_52),
    .io_validout64_53(middle_io_validout64_53),
    .io_validout64_54(middle_io_validout64_54),
    .io_validout64_55(middle_io_validout64_55),
    .io_validout64_56(middle_io_validout64_56),
    .io_validout64_57(middle_io_validout64_57),
    .io_validout64_58(middle_io_validout64_58),
    .io_validout64_59(middle_io_validout64_59),
    .io_validout64_60(middle_io_validout64_60),
    .io_validout64_61(middle_io_validout64_61),
    .io_validout64_62(middle_io_validout64_62),
    .io_validout64_63(middle_io_validout64_63),
    .io_tagout_Tag(middle_io_tagout_Tag),
    .io_tagout_RoundCnt(middle_io_tagout_RoundCnt),
    .io_addrout(middle_io_addrout),
    .io_ctrl(middle_io_ctrl)
  );
  CLOSegress1 egress1 ( // @[BuildingBlockNew.scala 87:23]
    .clock(egress1_clock),
    .io_in64_0(egress1_io_in64_0),
    .io_in64_1(egress1_io_in64_1),
    .io_in64_2(egress1_io_in64_2),
    .io_in64_3(egress1_io_in64_3),
    .io_in64_4(egress1_io_in64_4),
    .io_in64_5(egress1_io_in64_5),
    .io_in64_6(egress1_io_in64_6),
    .io_in64_7(egress1_io_in64_7),
    .io_in64_8(egress1_io_in64_8),
    .io_in64_9(egress1_io_in64_9),
    .io_in64_10(egress1_io_in64_10),
    .io_in64_11(egress1_io_in64_11),
    .io_in64_12(egress1_io_in64_12),
    .io_in64_13(egress1_io_in64_13),
    .io_in64_14(egress1_io_in64_14),
    .io_in64_15(egress1_io_in64_15),
    .io_in64_16(egress1_io_in64_16),
    .io_in64_17(egress1_io_in64_17),
    .io_in64_18(egress1_io_in64_18),
    .io_in64_19(egress1_io_in64_19),
    .io_in64_20(egress1_io_in64_20),
    .io_in64_21(egress1_io_in64_21),
    .io_in64_22(egress1_io_in64_22),
    .io_in64_23(egress1_io_in64_23),
    .io_in64_24(egress1_io_in64_24),
    .io_in64_25(egress1_io_in64_25),
    .io_in64_26(egress1_io_in64_26),
    .io_in64_27(egress1_io_in64_27),
    .io_in64_28(egress1_io_in64_28),
    .io_in64_29(egress1_io_in64_29),
    .io_in64_30(egress1_io_in64_30),
    .io_in64_31(egress1_io_in64_31),
    .io_in64_32(egress1_io_in64_32),
    .io_in64_33(egress1_io_in64_33),
    .io_in64_34(egress1_io_in64_34),
    .io_in64_35(egress1_io_in64_35),
    .io_in64_36(egress1_io_in64_36),
    .io_in64_37(egress1_io_in64_37),
    .io_in64_38(egress1_io_in64_38),
    .io_in64_39(egress1_io_in64_39),
    .io_in64_40(egress1_io_in64_40),
    .io_in64_41(egress1_io_in64_41),
    .io_in64_42(egress1_io_in64_42),
    .io_in64_43(egress1_io_in64_43),
    .io_in64_44(egress1_io_in64_44),
    .io_in64_45(egress1_io_in64_45),
    .io_in64_46(egress1_io_in64_46),
    .io_in64_47(egress1_io_in64_47),
    .io_in64_48(egress1_io_in64_48),
    .io_in64_49(egress1_io_in64_49),
    .io_in64_50(egress1_io_in64_50),
    .io_in64_51(egress1_io_in64_51),
    .io_in64_52(egress1_io_in64_52),
    .io_in64_53(egress1_io_in64_53),
    .io_in64_54(egress1_io_in64_54),
    .io_in64_55(egress1_io_in64_55),
    .io_in64_56(egress1_io_in64_56),
    .io_in64_57(egress1_io_in64_57),
    .io_in64_58(egress1_io_in64_58),
    .io_in64_59(egress1_io_in64_59),
    .io_in64_60(egress1_io_in64_60),
    .io_in64_61(egress1_io_in64_61),
    .io_in64_62(egress1_io_in64_62),
    .io_in64_63(egress1_io_in64_63),
    .io_validin64_0(egress1_io_validin64_0),
    .io_validin64_1(egress1_io_validin64_1),
    .io_validin64_2(egress1_io_validin64_2),
    .io_validin64_3(egress1_io_validin64_3),
    .io_validin64_4(egress1_io_validin64_4),
    .io_validin64_5(egress1_io_validin64_5),
    .io_validin64_6(egress1_io_validin64_6),
    .io_validin64_7(egress1_io_validin64_7),
    .io_validin64_8(egress1_io_validin64_8),
    .io_validin64_9(egress1_io_validin64_9),
    .io_validin64_10(egress1_io_validin64_10),
    .io_validin64_11(egress1_io_validin64_11),
    .io_validin64_12(egress1_io_validin64_12),
    .io_validin64_13(egress1_io_validin64_13),
    .io_validin64_14(egress1_io_validin64_14),
    .io_validin64_15(egress1_io_validin64_15),
    .io_validin64_16(egress1_io_validin64_16),
    .io_validin64_17(egress1_io_validin64_17),
    .io_validin64_18(egress1_io_validin64_18),
    .io_validin64_19(egress1_io_validin64_19),
    .io_validin64_20(egress1_io_validin64_20),
    .io_validin64_21(egress1_io_validin64_21),
    .io_validin64_22(egress1_io_validin64_22),
    .io_validin64_23(egress1_io_validin64_23),
    .io_validin64_24(egress1_io_validin64_24),
    .io_validin64_25(egress1_io_validin64_25),
    .io_validin64_26(egress1_io_validin64_26),
    .io_validin64_27(egress1_io_validin64_27),
    .io_validin64_28(egress1_io_validin64_28),
    .io_validin64_29(egress1_io_validin64_29),
    .io_validin64_30(egress1_io_validin64_30),
    .io_validin64_31(egress1_io_validin64_31),
    .io_validin64_32(egress1_io_validin64_32),
    .io_validin64_33(egress1_io_validin64_33),
    .io_validin64_34(egress1_io_validin64_34),
    .io_validin64_35(egress1_io_validin64_35),
    .io_validin64_36(egress1_io_validin64_36),
    .io_validin64_37(egress1_io_validin64_37),
    .io_validin64_38(egress1_io_validin64_38),
    .io_validin64_39(egress1_io_validin64_39),
    .io_validin64_40(egress1_io_validin64_40),
    .io_validin64_41(egress1_io_validin64_41),
    .io_validin64_42(egress1_io_validin64_42),
    .io_validin64_43(egress1_io_validin64_43),
    .io_validin64_44(egress1_io_validin64_44),
    .io_validin64_45(egress1_io_validin64_45),
    .io_validin64_46(egress1_io_validin64_46),
    .io_validin64_47(egress1_io_validin64_47),
    .io_validin64_48(egress1_io_validin64_48),
    .io_validin64_49(egress1_io_validin64_49),
    .io_validin64_50(egress1_io_validin64_50),
    .io_validin64_51(egress1_io_validin64_51),
    .io_validin64_52(egress1_io_validin64_52),
    .io_validin64_53(egress1_io_validin64_53),
    .io_validin64_54(egress1_io_validin64_54),
    .io_validin64_55(egress1_io_validin64_55),
    .io_validin64_56(egress1_io_validin64_56),
    .io_validin64_57(egress1_io_validin64_57),
    .io_validin64_58(egress1_io_validin64_58),
    .io_validin64_59(egress1_io_validin64_59),
    .io_validin64_60(egress1_io_validin64_60),
    .io_validin64_61(egress1_io_validin64_61),
    .io_validin64_62(egress1_io_validin64_62),
    .io_validin64_63(egress1_io_validin64_63),
    .io_tagin_Tag(egress1_io_tagin_Tag),
    .io_tagin_RoundCnt(egress1_io_tagin_RoundCnt),
    .io_addrin(egress1_io_addrin),
    .io_out64_0(egress1_io_out64_0),
    .io_out64_1(egress1_io_out64_1),
    .io_out64_2(egress1_io_out64_2),
    .io_out64_3(egress1_io_out64_3),
    .io_out64_4(egress1_io_out64_4),
    .io_out64_5(egress1_io_out64_5),
    .io_out64_6(egress1_io_out64_6),
    .io_out64_7(egress1_io_out64_7),
    .io_out64_8(egress1_io_out64_8),
    .io_out64_9(egress1_io_out64_9),
    .io_out64_10(egress1_io_out64_10),
    .io_out64_11(egress1_io_out64_11),
    .io_out64_12(egress1_io_out64_12),
    .io_out64_13(egress1_io_out64_13),
    .io_out64_14(egress1_io_out64_14),
    .io_out64_15(egress1_io_out64_15),
    .io_out64_16(egress1_io_out64_16),
    .io_out64_17(egress1_io_out64_17),
    .io_out64_18(egress1_io_out64_18),
    .io_out64_19(egress1_io_out64_19),
    .io_out64_20(egress1_io_out64_20),
    .io_out64_21(egress1_io_out64_21),
    .io_out64_22(egress1_io_out64_22),
    .io_out64_23(egress1_io_out64_23),
    .io_out64_24(egress1_io_out64_24),
    .io_out64_25(egress1_io_out64_25),
    .io_out64_26(egress1_io_out64_26),
    .io_out64_27(egress1_io_out64_27),
    .io_out64_28(egress1_io_out64_28),
    .io_out64_29(egress1_io_out64_29),
    .io_out64_30(egress1_io_out64_30),
    .io_out64_31(egress1_io_out64_31),
    .io_out64_32(egress1_io_out64_32),
    .io_out64_33(egress1_io_out64_33),
    .io_out64_34(egress1_io_out64_34),
    .io_out64_35(egress1_io_out64_35),
    .io_out64_36(egress1_io_out64_36),
    .io_out64_37(egress1_io_out64_37),
    .io_out64_38(egress1_io_out64_38),
    .io_out64_39(egress1_io_out64_39),
    .io_out64_40(egress1_io_out64_40),
    .io_out64_41(egress1_io_out64_41),
    .io_out64_42(egress1_io_out64_42),
    .io_out64_43(egress1_io_out64_43),
    .io_out64_44(egress1_io_out64_44),
    .io_out64_45(egress1_io_out64_45),
    .io_out64_46(egress1_io_out64_46),
    .io_out64_47(egress1_io_out64_47),
    .io_out64_48(egress1_io_out64_48),
    .io_out64_49(egress1_io_out64_49),
    .io_out64_50(egress1_io_out64_50),
    .io_out64_51(egress1_io_out64_51),
    .io_out64_52(egress1_io_out64_52),
    .io_out64_53(egress1_io_out64_53),
    .io_out64_54(egress1_io_out64_54),
    .io_out64_55(egress1_io_out64_55),
    .io_out64_56(egress1_io_out64_56),
    .io_out64_57(egress1_io_out64_57),
    .io_out64_58(egress1_io_out64_58),
    .io_out64_59(egress1_io_out64_59),
    .io_out64_60(egress1_io_out64_60),
    .io_out64_61(egress1_io_out64_61),
    .io_out64_62(egress1_io_out64_62),
    .io_out64_63(egress1_io_out64_63),
    .io_validout64_0(egress1_io_validout64_0),
    .io_validout64_1(egress1_io_validout64_1),
    .io_validout64_2(egress1_io_validout64_2),
    .io_validout64_3(egress1_io_validout64_3),
    .io_validout64_4(egress1_io_validout64_4),
    .io_validout64_5(egress1_io_validout64_5),
    .io_validout64_6(egress1_io_validout64_6),
    .io_validout64_7(egress1_io_validout64_7),
    .io_validout64_8(egress1_io_validout64_8),
    .io_validout64_9(egress1_io_validout64_9),
    .io_validout64_10(egress1_io_validout64_10),
    .io_validout64_11(egress1_io_validout64_11),
    .io_validout64_12(egress1_io_validout64_12),
    .io_validout64_13(egress1_io_validout64_13),
    .io_validout64_14(egress1_io_validout64_14),
    .io_validout64_15(egress1_io_validout64_15),
    .io_validout64_16(egress1_io_validout64_16),
    .io_validout64_17(egress1_io_validout64_17),
    .io_validout64_18(egress1_io_validout64_18),
    .io_validout64_19(egress1_io_validout64_19),
    .io_validout64_20(egress1_io_validout64_20),
    .io_validout64_21(egress1_io_validout64_21),
    .io_validout64_22(egress1_io_validout64_22),
    .io_validout64_23(egress1_io_validout64_23),
    .io_validout64_24(egress1_io_validout64_24),
    .io_validout64_25(egress1_io_validout64_25),
    .io_validout64_26(egress1_io_validout64_26),
    .io_validout64_27(egress1_io_validout64_27),
    .io_validout64_28(egress1_io_validout64_28),
    .io_validout64_29(egress1_io_validout64_29),
    .io_validout64_30(egress1_io_validout64_30),
    .io_validout64_31(egress1_io_validout64_31),
    .io_validout64_32(egress1_io_validout64_32),
    .io_validout64_33(egress1_io_validout64_33),
    .io_validout64_34(egress1_io_validout64_34),
    .io_validout64_35(egress1_io_validout64_35),
    .io_validout64_36(egress1_io_validout64_36),
    .io_validout64_37(egress1_io_validout64_37),
    .io_validout64_38(egress1_io_validout64_38),
    .io_validout64_39(egress1_io_validout64_39),
    .io_validout64_40(egress1_io_validout64_40),
    .io_validout64_41(egress1_io_validout64_41),
    .io_validout64_42(egress1_io_validout64_42),
    .io_validout64_43(egress1_io_validout64_43),
    .io_validout64_44(egress1_io_validout64_44),
    .io_validout64_45(egress1_io_validout64_45),
    .io_validout64_46(egress1_io_validout64_46),
    .io_validout64_47(egress1_io_validout64_47),
    .io_validout64_48(egress1_io_validout64_48),
    .io_validout64_49(egress1_io_validout64_49),
    .io_validout64_50(egress1_io_validout64_50),
    .io_validout64_51(egress1_io_validout64_51),
    .io_validout64_52(egress1_io_validout64_52),
    .io_validout64_53(egress1_io_validout64_53),
    .io_validout64_54(egress1_io_validout64_54),
    .io_validout64_55(egress1_io_validout64_55),
    .io_validout64_56(egress1_io_validout64_56),
    .io_validout64_57(egress1_io_validout64_57),
    .io_validout64_58(egress1_io_validout64_58),
    .io_validout64_59(egress1_io_validout64_59),
    .io_validout64_60(egress1_io_validout64_60),
    .io_validout64_61(egress1_io_validout64_61),
    .io_validout64_62(egress1_io_validout64_62),
    .io_validout64_63(egress1_io_validout64_63),
    .io_tagout_Tag(egress1_io_tagout_Tag),
    .io_tagout_RoundCnt(egress1_io_tagout_RoundCnt),
    .io_addrout(egress1_io_addrout),
    .io_ctrl(egress1_io_ctrl)
  );
  CLOSegress2 egress2 ( // @[BuildingBlockNew.scala 88:23]
    .clock(egress2_clock),
    .io_in64_0(egress2_io_in64_0),
    .io_in64_1(egress2_io_in64_1),
    .io_in64_2(egress2_io_in64_2),
    .io_in64_3(egress2_io_in64_3),
    .io_in64_4(egress2_io_in64_4),
    .io_in64_5(egress2_io_in64_5),
    .io_in64_6(egress2_io_in64_6),
    .io_in64_7(egress2_io_in64_7),
    .io_in64_8(egress2_io_in64_8),
    .io_in64_9(egress2_io_in64_9),
    .io_in64_10(egress2_io_in64_10),
    .io_in64_11(egress2_io_in64_11),
    .io_in64_12(egress2_io_in64_12),
    .io_in64_13(egress2_io_in64_13),
    .io_in64_14(egress2_io_in64_14),
    .io_in64_15(egress2_io_in64_15),
    .io_in64_16(egress2_io_in64_16),
    .io_in64_17(egress2_io_in64_17),
    .io_in64_18(egress2_io_in64_18),
    .io_in64_19(egress2_io_in64_19),
    .io_in64_20(egress2_io_in64_20),
    .io_in64_21(egress2_io_in64_21),
    .io_in64_22(egress2_io_in64_22),
    .io_in64_23(egress2_io_in64_23),
    .io_in64_24(egress2_io_in64_24),
    .io_in64_25(egress2_io_in64_25),
    .io_in64_26(egress2_io_in64_26),
    .io_in64_27(egress2_io_in64_27),
    .io_in64_28(egress2_io_in64_28),
    .io_in64_29(egress2_io_in64_29),
    .io_in64_30(egress2_io_in64_30),
    .io_in64_31(egress2_io_in64_31),
    .io_in64_32(egress2_io_in64_32),
    .io_in64_33(egress2_io_in64_33),
    .io_in64_34(egress2_io_in64_34),
    .io_in64_35(egress2_io_in64_35),
    .io_in64_36(egress2_io_in64_36),
    .io_in64_37(egress2_io_in64_37),
    .io_in64_38(egress2_io_in64_38),
    .io_in64_39(egress2_io_in64_39),
    .io_in64_40(egress2_io_in64_40),
    .io_in64_41(egress2_io_in64_41),
    .io_in64_42(egress2_io_in64_42),
    .io_in64_43(egress2_io_in64_43),
    .io_in64_44(egress2_io_in64_44),
    .io_in64_45(egress2_io_in64_45),
    .io_in64_46(egress2_io_in64_46),
    .io_in64_47(egress2_io_in64_47),
    .io_in64_48(egress2_io_in64_48),
    .io_in64_49(egress2_io_in64_49),
    .io_in64_50(egress2_io_in64_50),
    .io_in64_51(egress2_io_in64_51),
    .io_in64_52(egress2_io_in64_52),
    .io_in64_53(egress2_io_in64_53),
    .io_in64_54(egress2_io_in64_54),
    .io_in64_55(egress2_io_in64_55),
    .io_in64_56(egress2_io_in64_56),
    .io_in64_57(egress2_io_in64_57),
    .io_in64_58(egress2_io_in64_58),
    .io_in64_59(egress2_io_in64_59),
    .io_in64_60(egress2_io_in64_60),
    .io_in64_61(egress2_io_in64_61),
    .io_in64_62(egress2_io_in64_62),
    .io_in64_63(egress2_io_in64_63),
    .io_validin64_0(egress2_io_validin64_0),
    .io_validin64_1(egress2_io_validin64_1),
    .io_validin64_2(egress2_io_validin64_2),
    .io_validin64_3(egress2_io_validin64_3),
    .io_validin64_4(egress2_io_validin64_4),
    .io_validin64_5(egress2_io_validin64_5),
    .io_validin64_6(egress2_io_validin64_6),
    .io_validin64_7(egress2_io_validin64_7),
    .io_validin64_8(egress2_io_validin64_8),
    .io_validin64_9(egress2_io_validin64_9),
    .io_validin64_10(egress2_io_validin64_10),
    .io_validin64_11(egress2_io_validin64_11),
    .io_validin64_12(egress2_io_validin64_12),
    .io_validin64_13(egress2_io_validin64_13),
    .io_validin64_14(egress2_io_validin64_14),
    .io_validin64_15(egress2_io_validin64_15),
    .io_validin64_16(egress2_io_validin64_16),
    .io_validin64_17(egress2_io_validin64_17),
    .io_validin64_18(egress2_io_validin64_18),
    .io_validin64_19(egress2_io_validin64_19),
    .io_validin64_20(egress2_io_validin64_20),
    .io_validin64_21(egress2_io_validin64_21),
    .io_validin64_22(egress2_io_validin64_22),
    .io_validin64_23(egress2_io_validin64_23),
    .io_validin64_24(egress2_io_validin64_24),
    .io_validin64_25(egress2_io_validin64_25),
    .io_validin64_26(egress2_io_validin64_26),
    .io_validin64_27(egress2_io_validin64_27),
    .io_validin64_28(egress2_io_validin64_28),
    .io_validin64_29(egress2_io_validin64_29),
    .io_validin64_30(egress2_io_validin64_30),
    .io_validin64_31(egress2_io_validin64_31),
    .io_validin64_32(egress2_io_validin64_32),
    .io_validin64_33(egress2_io_validin64_33),
    .io_validin64_34(egress2_io_validin64_34),
    .io_validin64_35(egress2_io_validin64_35),
    .io_validin64_36(egress2_io_validin64_36),
    .io_validin64_37(egress2_io_validin64_37),
    .io_validin64_38(egress2_io_validin64_38),
    .io_validin64_39(egress2_io_validin64_39),
    .io_validin64_40(egress2_io_validin64_40),
    .io_validin64_41(egress2_io_validin64_41),
    .io_validin64_42(egress2_io_validin64_42),
    .io_validin64_43(egress2_io_validin64_43),
    .io_validin64_44(egress2_io_validin64_44),
    .io_validin64_45(egress2_io_validin64_45),
    .io_validin64_46(egress2_io_validin64_46),
    .io_validin64_47(egress2_io_validin64_47),
    .io_validin64_48(egress2_io_validin64_48),
    .io_validin64_49(egress2_io_validin64_49),
    .io_validin64_50(egress2_io_validin64_50),
    .io_validin64_51(egress2_io_validin64_51),
    .io_validin64_52(egress2_io_validin64_52),
    .io_validin64_53(egress2_io_validin64_53),
    .io_validin64_54(egress2_io_validin64_54),
    .io_validin64_55(egress2_io_validin64_55),
    .io_validin64_56(egress2_io_validin64_56),
    .io_validin64_57(egress2_io_validin64_57),
    .io_validin64_58(egress2_io_validin64_58),
    .io_validin64_59(egress2_io_validin64_59),
    .io_validin64_60(egress2_io_validin64_60),
    .io_validin64_61(egress2_io_validin64_61),
    .io_validin64_62(egress2_io_validin64_62),
    .io_validin64_63(egress2_io_validin64_63),
    .io_tagin_Tag(egress2_io_tagin_Tag),
    .io_tagin_RoundCnt(egress2_io_tagin_RoundCnt),
    .io_addrin(egress2_io_addrin),
    .io_out64_0(egress2_io_out64_0),
    .io_out64_1(egress2_io_out64_1),
    .io_out64_2(egress2_io_out64_2),
    .io_out64_3(egress2_io_out64_3),
    .io_out64_4(egress2_io_out64_4),
    .io_out64_5(egress2_io_out64_5),
    .io_out64_6(egress2_io_out64_6),
    .io_out64_7(egress2_io_out64_7),
    .io_out64_8(egress2_io_out64_8),
    .io_out64_9(egress2_io_out64_9),
    .io_out64_10(egress2_io_out64_10),
    .io_out64_11(egress2_io_out64_11),
    .io_out64_12(egress2_io_out64_12),
    .io_out64_13(egress2_io_out64_13),
    .io_out64_14(egress2_io_out64_14),
    .io_out64_15(egress2_io_out64_15),
    .io_out64_16(egress2_io_out64_16),
    .io_out64_17(egress2_io_out64_17),
    .io_out64_18(egress2_io_out64_18),
    .io_out64_19(egress2_io_out64_19),
    .io_out64_20(egress2_io_out64_20),
    .io_out64_21(egress2_io_out64_21),
    .io_out64_22(egress2_io_out64_22),
    .io_out64_23(egress2_io_out64_23),
    .io_out64_24(egress2_io_out64_24),
    .io_out64_25(egress2_io_out64_25),
    .io_out64_26(egress2_io_out64_26),
    .io_out64_27(egress2_io_out64_27),
    .io_out64_28(egress2_io_out64_28),
    .io_out64_29(egress2_io_out64_29),
    .io_out64_30(egress2_io_out64_30),
    .io_out64_31(egress2_io_out64_31),
    .io_out64_32(egress2_io_out64_32),
    .io_out64_33(egress2_io_out64_33),
    .io_out64_34(egress2_io_out64_34),
    .io_out64_35(egress2_io_out64_35),
    .io_out64_36(egress2_io_out64_36),
    .io_out64_37(egress2_io_out64_37),
    .io_out64_38(egress2_io_out64_38),
    .io_out64_39(egress2_io_out64_39),
    .io_out64_40(egress2_io_out64_40),
    .io_out64_41(egress2_io_out64_41),
    .io_out64_42(egress2_io_out64_42),
    .io_out64_43(egress2_io_out64_43),
    .io_out64_44(egress2_io_out64_44),
    .io_out64_45(egress2_io_out64_45),
    .io_out64_46(egress2_io_out64_46),
    .io_out64_47(egress2_io_out64_47),
    .io_out64_48(egress2_io_out64_48),
    .io_out64_49(egress2_io_out64_49),
    .io_out64_50(egress2_io_out64_50),
    .io_out64_51(egress2_io_out64_51),
    .io_out64_52(egress2_io_out64_52),
    .io_out64_53(egress2_io_out64_53),
    .io_out64_54(egress2_io_out64_54),
    .io_out64_55(egress2_io_out64_55),
    .io_out64_56(egress2_io_out64_56),
    .io_out64_57(egress2_io_out64_57),
    .io_out64_58(egress2_io_out64_58),
    .io_out64_59(egress2_io_out64_59),
    .io_out64_60(egress2_io_out64_60),
    .io_out64_61(egress2_io_out64_61),
    .io_out64_62(egress2_io_out64_62),
    .io_out64_63(egress2_io_out64_63),
    .io_validout64_0(egress2_io_validout64_0),
    .io_validout64_1(egress2_io_validout64_1),
    .io_validout64_2(egress2_io_validout64_2),
    .io_validout64_3(egress2_io_validout64_3),
    .io_validout64_4(egress2_io_validout64_4),
    .io_validout64_5(egress2_io_validout64_5),
    .io_validout64_6(egress2_io_validout64_6),
    .io_validout64_7(egress2_io_validout64_7),
    .io_validout64_8(egress2_io_validout64_8),
    .io_validout64_9(egress2_io_validout64_9),
    .io_validout64_10(egress2_io_validout64_10),
    .io_validout64_11(egress2_io_validout64_11),
    .io_validout64_12(egress2_io_validout64_12),
    .io_validout64_13(egress2_io_validout64_13),
    .io_validout64_14(egress2_io_validout64_14),
    .io_validout64_15(egress2_io_validout64_15),
    .io_validout64_16(egress2_io_validout64_16),
    .io_validout64_17(egress2_io_validout64_17),
    .io_validout64_18(egress2_io_validout64_18),
    .io_validout64_19(egress2_io_validout64_19),
    .io_validout64_20(egress2_io_validout64_20),
    .io_validout64_21(egress2_io_validout64_21),
    .io_validout64_22(egress2_io_validout64_22),
    .io_validout64_23(egress2_io_validout64_23),
    .io_validout64_24(egress2_io_validout64_24),
    .io_validout64_25(egress2_io_validout64_25),
    .io_validout64_26(egress2_io_validout64_26),
    .io_validout64_27(egress2_io_validout64_27),
    .io_validout64_28(egress2_io_validout64_28),
    .io_validout64_29(egress2_io_validout64_29),
    .io_validout64_30(egress2_io_validout64_30),
    .io_validout64_31(egress2_io_validout64_31),
    .io_validout64_32(egress2_io_validout64_32),
    .io_validout64_33(egress2_io_validout64_33),
    .io_validout64_34(egress2_io_validout64_34),
    .io_validout64_35(egress2_io_validout64_35),
    .io_validout64_36(egress2_io_validout64_36),
    .io_validout64_37(egress2_io_validout64_37),
    .io_validout64_38(egress2_io_validout64_38),
    .io_validout64_39(egress2_io_validout64_39),
    .io_validout64_40(egress2_io_validout64_40),
    .io_validout64_41(egress2_io_validout64_41),
    .io_validout64_42(egress2_io_validout64_42),
    .io_validout64_43(egress2_io_validout64_43),
    .io_validout64_44(egress2_io_validout64_44),
    .io_validout64_45(egress2_io_validout64_45),
    .io_validout64_46(egress2_io_validout64_46),
    .io_validout64_47(egress2_io_validout64_47),
    .io_validout64_48(egress2_io_validout64_48),
    .io_validout64_49(egress2_io_validout64_49),
    .io_validout64_50(egress2_io_validout64_50),
    .io_validout64_51(egress2_io_validout64_51),
    .io_validout64_52(egress2_io_validout64_52),
    .io_validout64_53(egress2_io_validout64_53),
    .io_validout64_54(egress2_io_validout64_54),
    .io_validout64_55(egress2_io_validout64_55),
    .io_validout64_56(egress2_io_validout64_56),
    .io_validout64_57(egress2_io_validout64_57),
    .io_validout64_58(egress2_io_validout64_58),
    .io_validout64_59(egress2_io_validout64_59),
    .io_validout64_60(egress2_io_validout64_60),
    .io_validout64_61(egress2_io_validout64_61),
    .io_validout64_62(egress2_io_validout64_62),
    .io_validout64_63(egress2_io_validout64_63),
    .io_tagout_Tag(egress2_io_tagout_Tag),
    .io_tagout_RoundCnt(egress2_io_tagout_RoundCnt),
    .io_addrout(egress2_io_addrout),
    .io_ctrl(egress2_io_ctrl)
  );
  assign io_d_out_0_a = egress2_io_out64_0; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_0_valid_a = egress2_io_validout64_0; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_0_b = egress2_io_out64_1; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_0_valid_b = egress2_io_validout64_1; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_1_a = egress2_io_out64_2; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_1_valid_a = egress2_io_validout64_2; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_1_b = egress2_io_out64_3; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_1_valid_b = egress2_io_validout64_3; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_2_a = egress2_io_out64_4; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_2_valid_a = egress2_io_validout64_4; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_2_b = egress2_io_out64_5; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_2_valid_b = egress2_io_validout64_5; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_3_a = egress2_io_out64_6; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_3_valid_a = egress2_io_validout64_6; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_3_b = egress2_io_out64_7; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_3_valid_b = egress2_io_validout64_7; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_4_a = egress2_io_out64_8; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_4_valid_a = egress2_io_validout64_8; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_4_b = egress2_io_out64_9; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_4_valid_b = egress2_io_validout64_9; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_5_a = egress2_io_out64_10; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_5_valid_a = egress2_io_validout64_10; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_5_b = egress2_io_out64_11; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_5_valid_b = egress2_io_validout64_11; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_6_a = egress2_io_out64_12; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_6_valid_a = egress2_io_validout64_12; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_6_b = egress2_io_out64_13; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_6_valid_b = egress2_io_validout64_13; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_7_a = egress2_io_out64_14; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_7_valid_a = egress2_io_validout64_14; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_7_b = egress2_io_out64_15; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_7_valid_b = egress2_io_validout64_15; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_8_a = egress2_io_out64_16; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_8_valid_a = egress2_io_validout64_16; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_8_b = egress2_io_out64_17; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_8_valid_b = egress2_io_validout64_17; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_9_a = egress2_io_out64_18; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_9_valid_a = egress2_io_validout64_18; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_9_b = egress2_io_out64_19; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_9_valid_b = egress2_io_validout64_19; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_10_a = egress2_io_out64_20; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_10_valid_a = egress2_io_validout64_20; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_10_b = egress2_io_out64_21; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_10_valid_b = egress2_io_validout64_21; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_11_a = egress2_io_out64_22; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_11_valid_a = egress2_io_validout64_22; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_11_b = egress2_io_out64_23; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_11_valid_b = egress2_io_validout64_23; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_12_a = egress2_io_out64_24; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_12_valid_a = egress2_io_validout64_24; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_12_b = egress2_io_out64_25; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_12_valid_b = egress2_io_validout64_25; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_13_a = egress2_io_out64_26; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_13_valid_a = egress2_io_validout64_26; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_13_b = egress2_io_out64_27; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_13_valid_b = egress2_io_validout64_27; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_14_a = egress2_io_out64_28; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_14_valid_a = egress2_io_validout64_28; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_14_b = egress2_io_out64_29; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_14_valid_b = egress2_io_validout64_29; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_15_a = egress2_io_out64_30; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_15_valid_a = egress2_io_validout64_30; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_15_b = egress2_io_out64_31; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_15_valid_b = egress2_io_validout64_31; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_16_a = egress2_io_out64_32; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_16_valid_a = egress2_io_validout64_32; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_16_b = egress2_io_out64_33; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_16_valid_b = egress2_io_validout64_33; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_17_a = egress2_io_out64_34; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_17_valid_a = egress2_io_validout64_34; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_17_b = egress2_io_out64_35; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_17_valid_b = egress2_io_validout64_35; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_18_a = egress2_io_out64_36; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_18_valid_a = egress2_io_validout64_36; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_18_b = egress2_io_out64_37; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_18_valid_b = egress2_io_validout64_37; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_19_a = egress2_io_out64_38; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_19_valid_a = egress2_io_validout64_38; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_19_b = egress2_io_out64_39; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_19_valid_b = egress2_io_validout64_39; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_20_a = egress2_io_out64_40; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_20_valid_a = egress2_io_validout64_40; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_20_b = egress2_io_out64_41; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_20_valid_b = egress2_io_validout64_41; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_21_a = egress2_io_out64_42; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_21_valid_a = egress2_io_validout64_42; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_21_b = egress2_io_out64_43; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_21_valid_b = egress2_io_validout64_43; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_22_a = egress2_io_out64_44; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_22_valid_a = egress2_io_validout64_44; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_22_b = egress2_io_out64_45; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_22_valid_b = egress2_io_validout64_45; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_23_a = egress2_io_out64_46; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_23_valid_a = egress2_io_validout64_46; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_23_b = egress2_io_out64_47; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_23_valid_b = egress2_io_validout64_47; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_24_a = egress2_io_out64_48; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_24_valid_a = egress2_io_validout64_48; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_24_b = egress2_io_out64_49; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_24_valid_b = egress2_io_validout64_49; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_25_a = egress2_io_out64_50; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_25_valid_a = egress2_io_validout64_50; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_25_b = egress2_io_out64_51; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_25_valid_b = egress2_io_validout64_51; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_26_a = egress2_io_out64_52; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_26_valid_a = egress2_io_validout64_52; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_26_b = egress2_io_out64_53; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_26_valid_b = egress2_io_validout64_53; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_27_a = egress2_io_out64_54; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_27_valid_a = egress2_io_validout64_54; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_27_b = egress2_io_out64_55; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_27_valid_b = egress2_io_validout64_55; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_28_a = egress2_io_out64_56; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_28_valid_a = egress2_io_validout64_56; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_28_b = egress2_io_out64_57; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_28_valid_b = egress2_io_validout64_57; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_29_a = egress2_io_out64_58; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_29_valid_a = egress2_io_validout64_58; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_29_b = egress2_io_out64_59; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_29_valid_b = egress2_io_validout64_59; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_30_a = egress2_io_out64_60; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_30_valid_a = egress2_io_validout64_60; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_30_b = egress2_io_out64_61; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_30_valid_b = egress2_io_validout64_61; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_31_a = egress2_io_out64_62; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_31_valid_a = egress2_io_validout64_62; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_31_b = egress2_io_out64_63; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_31_valid_b = egress2_io_validout64_63; // @[BuildingBlockNew.scala 316:25]
  assign io_PC6_out = PC6; // @[BuildingBlockNew.scala 161:14]
  assign io_Addr_out = egress2_io_addrout; // @[BuildingBlockNew.scala 319:15]
  assign io_Tag_out_Tag = egress2_io_tagout_Tag; // @[BuildingBlockNew.scala 318:14]
  assign io_Tag_out_RoundCnt = egress2_io_tagout_RoundCnt; // @[BuildingBlockNew.scala 318:14]
  assign Mem1_R0_addr = io_wr_en_mem1 ? wrAddr1 : PC1; // @[BuildingBlockNew.scala 223:22 BuildingBlockNew.scala 225:14 BuildingBlockNew.scala 230:14]
  assign Mem1_R0_clk = clock; // @[BuildingBlockNew.scala 223:22 BuildingBlockNew.scala 229:24]
  assign Mem1_W0_addr = io_wr_en_mem1 ? wrAddr1 : PC1; // @[BuildingBlockNew.scala 223:22 BuildingBlockNew.scala 225:14 BuildingBlockNew.scala 230:14]
  assign Mem1_W0_en = io_wr_en_mem1; // @[BuildingBlockNew.scala 223:22 BuildingBlockNew.scala 34:25]
  assign Mem1_W0_clk = clock; // @[BuildingBlockNew.scala 223:22]
  assign Mem1_W0_data = io_wr_instr_mem1; // @[BuildingBlockNew.scala 223:22]
  assign Mem2_R0_addr = io_wr_en_mem2 ? wrAddr2 : PC2; // @[BuildingBlockNew.scala 232:22 BuildingBlockNew.scala 234:14 BuildingBlockNew.scala 239:14]
  assign Mem2_R0_clk = clock; // @[BuildingBlockNew.scala 232:22 BuildingBlockNew.scala 238:24]
  assign Mem2_W0_addr = io_wr_en_mem2 ? wrAddr2 : PC2; // @[BuildingBlockNew.scala 232:22 BuildingBlockNew.scala 234:14 BuildingBlockNew.scala 239:14]
  assign Mem2_W0_en = io_wr_en_mem2; // @[BuildingBlockNew.scala 232:22 BuildingBlockNew.scala 35:25]
  assign Mem2_W0_clk = clock; // @[BuildingBlockNew.scala 232:22]
  assign Mem2_W0_data = io_wr_instr_mem2; // @[BuildingBlockNew.scala 232:22]
  assign Mem3_R0_addr = io_wr_en_mem3 ? wrAddr3 : PC3; // @[BuildingBlockNew.scala 241:22 BuildingBlockNew.scala 243:14 BuildingBlockNew.scala 248:14]
  assign Mem3_R0_clk = clock; // @[BuildingBlockNew.scala 241:22 BuildingBlockNew.scala 247:24]
  assign Mem3_W0_addr = io_wr_en_mem3 ? wrAddr3 : PC3; // @[BuildingBlockNew.scala 241:22 BuildingBlockNew.scala 243:14 BuildingBlockNew.scala 248:14]
  assign Mem3_W0_en = io_wr_en_mem3; // @[BuildingBlockNew.scala 241:22 BuildingBlockNew.scala 36:25]
  assign Mem3_W0_clk = clock; // @[BuildingBlockNew.scala 241:22]
  assign Mem3_W0_data = io_wr_instr_mem3; // @[BuildingBlockNew.scala 241:22]
  assign Mem4_R0_addr = io_wr_en_mem4 ? wrAddr4 : PC4; // @[BuildingBlockNew.scala 250:22 BuildingBlockNew.scala 252:14 BuildingBlockNew.scala 257:14]
  assign Mem4_R0_clk = clock; // @[BuildingBlockNew.scala 250:22 BuildingBlockNew.scala 256:24]
  assign Mem4_W0_addr = io_wr_en_mem4 ? wrAddr4 : PC4; // @[BuildingBlockNew.scala 250:22 BuildingBlockNew.scala 252:14 BuildingBlockNew.scala 257:14]
  assign Mem4_W0_en = io_wr_en_mem4; // @[BuildingBlockNew.scala 250:22 BuildingBlockNew.scala 37:25]
  assign Mem4_W0_clk = clock; // @[BuildingBlockNew.scala 250:22]
  assign Mem4_W0_data = io_wr_instr_mem4; // @[BuildingBlockNew.scala 250:22]
  assign Mem5_R0_addr = io_wr_en_mem5 ? wrAddr5 : PC5; // @[BuildingBlockNew.scala 259:22 BuildingBlockNew.scala 261:14 BuildingBlockNew.scala 266:14]
  assign Mem5_R0_clk = clock; // @[BuildingBlockNew.scala 259:22 BuildingBlockNew.scala 265:24]
  assign Mem5_W0_addr = io_wr_en_mem5 ? wrAddr5 : PC5; // @[BuildingBlockNew.scala 259:22 BuildingBlockNew.scala 261:14 BuildingBlockNew.scala 266:14]
  assign Mem5_W0_en = io_wr_en_mem5; // @[BuildingBlockNew.scala 259:22 BuildingBlockNew.scala 38:25]
  assign Mem5_W0_clk = clock; // @[BuildingBlockNew.scala 259:22]
  assign Mem5_W0_data = io_wr_instr_mem5; // @[BuildingBlockNew.scala 259:22]
  assign Mem6_R0_addr = io_wr_en_mem6 ? wrAddr6 : PC6; // @[BuildingBlockNew.scala 268:22 BuildingBlockNew.scala 270:14 BuildingBlockNew.scala 275:14]
  assign Mem6_R0_clk = clock; // @[BuildingBlockNew.scala 268:22 BuildingBlockNew.scala 274:24]
  assign Mem6_W0_addr = io_wr_en_mem6 ? wrAddr6 : PC6; // @[BuildingBlockNew.scala 268:22 BuildingBlockNew.scala 270:14 BuildingBlockNew.scala 275:14]
  assign Mem6_W0_en = io_wr_en_mem6; // @[BuildingBlockNew.scala 268:22 BuildingBlockNew.scala 39:25]
  assign Mem6_W0_clk = clock; // @[BuildingBlockNew.scala 268:22]
  assign Mem6_W0_data = io_wr_instr_mem6; // @[BuildingBlockNew.scala 268:22]
  assign peCol_clock = clock;
  assign peCol_reset = reset;
  assign peCol_io_d_in_0_a = io_d_in_0_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_0_valid_a = io_d_in_0_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_0_b = io_d_in_0_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_1_a = io_d_in_1_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_1_valid_a = io_d_in_1_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_1_b = io_d_in_1_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_2_a = io_d_in_2_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_2_valid_a = io_d_in_2_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_2_b = io_d_in_2_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_3_a = io_d_in_3_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_3_valid_a = io_d_in_3_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_3_b = io_d_in_3_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_4_a = io_d_in_4_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_4_valid_a = io_d_in_4_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_4_b = io_d_in_4_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_5_a = io_d_in_5_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_5_valid_a = io_d_in_5_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_5_b = io_d_in_5_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_6_a = io_d_in_6_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_6_valid_a = io_d_in_6_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_6_b = io_d_in_6_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_7_a = io_d_in_7_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_7_valid_a = io_d_in_7_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_7_b = io_d_in_7_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_8_a = io_d_in_8_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_8_valid_a = io_d_in_8_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_8_b = io_d_in_8_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_9_a = io_d_in_9_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_9_valid_a = io_d_in_9_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_9_b = io_d_in_9_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_10_a = io_d_in_10_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_10_valid_a = io_d_in_10_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_10_b = io_d_in_10_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_11_a = io_d_in_11_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_11_valid_a = io_d_in_11_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_11_b = io_d_in_11_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_12_a = io_d_in_12_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_12_valid_a = io_d_in_12_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_12_b = io_d_in_12_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_13_a = io_d_in_13_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_13_valid_a = io_d_in_13_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_13_b = io_d_in_13_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_14_a = io_d_in_14_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_14_valid_a = io_d_in_14_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_14_b = io_d_in_14_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_15_a = io_d_in_15_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_15_valid_a = io_d_in_15_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_15_b = io_d_in_15_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_16_a = io_d_in_16_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_16_valid_a = io_d_in_16_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_16_b = io_d_in_16_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_17_a = io_d_in_17_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_17_valid_a = io_d_in_17_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_17_b = io_d_in_17_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_18_a = io_d_in_18_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_18_valid_a = io_d_in_18_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_18_b = io_d_in_18_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_19_a = io_d_in_19_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_19_valid_a = io_d_in_19_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_19_b = io_d_in_19_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_20_a = io_d_in_20_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_20_valid_a = io_d_in_20_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_20_b = io_d_in_20_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_21_a = io_d_in_21_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_21_valid_a = io_d_in_21_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_21_b = io_d_in_21_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_22_a = io_d_in_22_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_22_valid_a = io_d_in_22_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_22_b = io_d_in_22_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_23_a = io_d_in_23_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_23_valid_a = io_d_in_23_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_23_b = io_d_in_23_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_24_a = io_d_in_24_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_24_valid_a = io_d_in_24_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_24_b = io_d_in_24_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_25_a = io_d_in_25_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_25_valid_a = io_d_in_25_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_25_b = io_d_in_25_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_26_a = io_d_in_26_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_26_valid_a = io_d_in_26_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_26_b = io_d_in_26_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_27_a = io_d_in_27_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_27_valid_a = io_d_in_27_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_27_b = io_d_in_27_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_28_a = io_d_in_28_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_28_valid_a = io_d_in_28_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_28_b = io_d_in_28_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_29_a = io_d_in_29_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_29_valid_a = io_d_in_29_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_29_b = io_d_in_29_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_30_a = io_d_in_30_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_30_valid_a = io_d_in_30_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_30_b = io_d_in_30_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_31_a = io_d_in_31_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_31_valid_a = io_d_in_31_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_31_b = io_d_in_31_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_tagin_Tag = io_Tag_in_Tag; // @[BuildingBlockNew.scala 281:18]
  assign peCol_io_tagin_RoundCnt = io_Tag_in_RoundCnt; // @[BuildingBlockNew.scala 281:18]
  assign peCol_io_addrin = io_Addr_in; // @[BuildingBlockNew.scala 282:19]
  assign peCol_io_instr = instr1; // @[BuildingBlockNew.scala 163:18]
  assign ingress1_clock = clock;
  assign ingress1_io_in64_0 = peCol_io_d_out_0_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_1 = peCol_io_d_out_0_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_2 = peCol_io_d_out_1_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_3 = peCol_io_d_out_1_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_4 = peCol_io_d_out_2_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_5 = peCol_io_d_out_2_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_6 = peCol_io_d_out_3_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_7 = peCol_io_d_out_3_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_8 = peCol_io_d_out_4_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_9 = peCol_io_d_out_4_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_10 = peCol_io_d_out_5_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_11 = peCol_io_d_out_5_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_12 = peCol_io_d_out_6_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_13 = peCol_io_d_out_6_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_14 = peCol_io_d_out_7_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_15 = peCol_io_d_out_7_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_16 = peCol_io_d_out_8_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_17 = peCol_io_d_out_8_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_18 = peCol_io_d_out_9_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_19 = peCol_io_d_out_9_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_20 = peCol_io_d_out_10_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_21 = peCol_io_d_out_10_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_22 = peCol_io_d_out_11_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_23 = peCol_io_d_out_11_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_24 = peCol_io_d_out_12_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_25 = peCol_io_d_out_12_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_26 = peCol_io_d_out_13_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_27 = peCol_io_d_out_13_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_28 = peCol_io_d_out_14_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_29 = peCol_io_d_out_14_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_30 = peCol_io_d_out_15_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_31 = peCol_io_d_out_15_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_32 = peCol_io_d_out_16_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_33 = peCol_io_d_out_16_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_34 = peCol_io_d_out_17_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_35 = peCol_io_d_out_17_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_36 = peCol_io_d_out_18_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_37 = peCol_io_d_out_18_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_38 = peCol_io_d_out_19_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_39 = peCol_io_d_out_19_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_40 = peCol_io_d_out_20_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_41 = peCol_io_d_out_20_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_42 = peCol_io_d_out_21_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_43 = peCol_io_d_out_21_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_44 = peCol_io_d_out_22_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_45 = peCol_io_d_out_22_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_46 = peCol_io_d_out_23_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_47 = peCol_io_d_out_23_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_48 = peCol_io_d_out_24_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_49 = peCol_io_d_out_24_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_50 = peCol_io_d_out_25_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_51 = peCol_io_d_out_25_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_52 = peCol_io_d_out_26_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_53 = peCol_io_d_out_26_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_54 = peCol_io_d_out_27_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_55 = peCol_io_d_out_27_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_56 = peCol_io_d_out_28_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_57 = peCol_io_d_out_28_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_58 = peCol_io_d_out_29_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_59 = peCol_io_d_out_29_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_60 = peCol_io_d_out_30_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_61 = peCol_io_d_out_30_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_62 = peCol_io_d_out_31_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_63 = peCol_io_d_out_31_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_validin64_0 = peCol_io_d_out_0_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_2 = peCol_io_d_out_1_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_4 = peCol_io_d_out_2_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_6 = peCol_io_d_out_3_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_8 = peCol_io_d_out_4_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_10 = peCol_io_d_out_5_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_12 = peCol_io_d_out_6_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_14 = peCol_io_d_out_7_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_16 = peCol_io_d_out_8_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_18 = peCol_io_d_out_9_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_20 = peCol_io_d_out_10_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_22 = peCol_io_d_out_11_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_24 = peCol_io_d_out_12_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_26 = peCol_io_d_out_13_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_28 = peCol_io_d_out_14_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_30 = peCol_io_d_out_15_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_32 = peCol_io_d_out_16_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_34 = peCol_io_d_out_17_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_36 = peCol_io_d_out_18_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_38 = peCol_io_d_out_19_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_40 = peCol_io_d_out_20_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_42 = peCol_io_d_out_21_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_44 = peCol_io_d_out_22_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_46 = peCol_io_d_out_23_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_48 = peCol_io_d_out_24_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_50 = peCol_io_d_out_25_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_52 = peCol_io_d_out_26_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_54 = peCol_io_d_out_27_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_56 = peCol_io_d_out_28_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_58 = peCol_io_d_out_29_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_60 = peCol_io_d_out_30_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_62 = peCol_io_d_out_31_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_tagin_Tag = peCol_io_tagout_Tag; // @[BuildingBlockNew.scala 284:21]
  assign ingress1_io_tagin_RoundCnt = peCol_io_tagout_RoundCnt; // @[BuildingBlockNew.scala 284:21]
  assign ingress1_io_addrin = peCol_io_addrout; // @[BuildingBlockNew.scala 285:22]
  assign ingress1_io_ctrl = instr2; // @[BuildingBlockNew.scala 164:20]
  assign ingress2_clock = clock;
  assign ingress2_io_in64_0 = ingress1_io_out64_0; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_1 = ingress1_io_out64_1; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_2 = ingress1_io_out64_2; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_3 = ingress1_io_out64_3; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_4 = ingress1_io_out64_4; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_5 = ingress1_io_out64_5; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_6 = ingress1_io_out64_6; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_7 = ingress1_io_out64_7; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_8 = ingress1_io_out64_8; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_9 = ingress1_io_out64_9; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_10 = ingress1_io_out64_10; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_11 = ingress1_io_out64_11; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_12 = ingress1_io_out64_12; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_13 = ingress1_io_out64_13; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_14 = ingress1_io_out64_14; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_15 = ingress1_io_out64_15; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_16 = ingress1_io_out64_16; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_17 = ingress1_io_out64_17; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_18 = ingress1_io_out64_18; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_19 = ingress1_io_out64_19; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_20 = ingress1_io_out64_20; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_21 = ingress1_io_out64_21; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_22 = ingress1_io_out64_22; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_23 = ingress1_io_out64_23; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_24 = ingress1_io_out64_24; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_25 = ingress1_io_out64_25; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_26 = ingress1_io_out64_26; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_27 = ingress1_io_out64_27; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_28 = ingress1_io_out64_28; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_29 = ingress1_io_out64_29; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_30 = ingress1_io_out64_30; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_31 = ingress1_io_out64_31; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_32 = ingress1_io_out64_32; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_33 = ingress1_io_out64_33; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_34 = ingress1_io_out64_34; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_35 = ingress1_io_out64_35; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_36 = ingress1_io_out64_36; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_37 = ingress1_io_out64_37; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_38 = ingress1_io_out64_38; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_39 = ingress1_io_out64_39; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_40 = ingress1_io_out64_40; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_41 = ingress1_io_out64_41; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_42 = ingress1_io_out64_42; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_43 = ingress1_io_out64_43; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_44 = ingress1_io_out64_44; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_45 = ingress1_io_out64_45; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_46 = ingress1_io_out64_46; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_47 = ingress1_io_out64_47; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_48 = ingress1_io_out64_48; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_49 = ingress1_io_out64_49; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_50 = ingress1_io_out64_50; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_51 = ingress1_io_out64_51; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_52 = ingress1_io_out64_52; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_53 = ingress1_io_out64_53; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_54 = ingress1_io_out64_54; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_55 = ingress1_io_out64_55; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_56 = ingress1_io_out64_56; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_57 = ingress1_io_out64_57; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_58 = ingress1_io_out64_58; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_59 = ingress1_io_out64_59; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_60 = ingress1_io_out64_60; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_61 = ingress1_io_out64_61; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_62 = ingress1_io_out64_62; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_63 = ingress1_io_out64_63; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_validin64_0 = ingress1_io_validout64_0; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_1 = ingress1_io_validout64_1; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_2 = ingress1_io_validout64_2; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_3 = ingress1_io_validout64_3; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_4 = ingress1_io_validout64_4; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_5 = ingress1_io_validout64_5; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_6 = ingress1_io_validout64_6; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_7 = ingress1_io_validout64_7; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_8 = ingress1_io_validout64_8; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_9 = ingress1_io_validout64_9; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_10 = ingress1_io_validout64_10; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_11 = ingress1_io_validout64_11; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_12 = ingress1_io_validout64_12; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_13 = ingress1_io_validout64_13; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_14 = ingress1_io_validout64_14; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_15 = ingress1_io_validout64_15; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_16 = ingress1_io_validout64_16; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_17 = ingress1_io_validout64_17; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_18 = ingress1_io_validout64_18; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_19 = ingress1_io_validout64_19; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_20 = ingress1_io_validout64_20; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_21 = ingress1_io_validout64_21; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_22 = ingress1_io_validout64_22; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_23 = ingress1_io_validout64_23; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_24 = ingress1_io_validout64_24; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_25 = ingress1_io_validout64_25; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_26 = ingress1_io_validout64_26; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_27 = ingress1_io_validout64_27; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_28 = ingress1_io_validout64_28; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_29 = ingress1_io_validout64_29; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_30 = ingress1_io_validout64_30; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_31 = ingress1_io_validout64_31; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_32 = ingress1_io_validout64_32; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_33 = ingress1_io_validout64_33; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_34 = ingress1_io_validout64_34; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_35 = ingress1_io_validout64_35; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_36 = ingress1_io_validout64_36; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_37 = ingress1_io_validout64_37; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_38 = ingress1_io_validout64_38; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_39 = ingress1_io_validout64_39; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_40 = ingress1_io_validout64_40; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_41 = ingress1_io_validout64_41; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_42 = ingress1_io_validout64_42; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_43 = ingress1_io_validout64_43; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_44 = ingress1_io_validout64_44; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_45 = ingress1_io_validout64_45; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_46 = ingress1_io_validout64_46; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_47 = ingress1_io_validout64_47; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_48 = ingress1_io_validout64_48; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_49 = ingress1_io_validout64_49; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_50 = ingress1_io_validout64_50; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_51 = ingress1_io_validout64_51; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_52 = ingress1_io_validout64_52; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_53 = ingress1_io_validout64_53; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_54 = ingress1_io_validout64_54; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_55 = ingress1_io_validout64_55; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_56 = ingress1_io_validout64_56; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_57 = ingress1_io_validout64_57; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_58 = ingress1_io_validout64_58; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_59 = ingress1_io_validout64_59; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_60 = ingress1_io_validout64_60; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_61 = ingress1_io_validout64_61; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_62 = ingress1_io_validout64_62; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_63 = ingress1_io_validout64_63; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_tagin_Tag = ingress1_io_tagout_Tag; // @[BuildingBlockNew.scala 295:21]
  assign ingress2_io_tagin_RoundCnt = ingress1_io_tagout_RoundCnt; // @[BuildingBlockNew.scala 295:21]
  assign ingress2_io_addrin = ingress1_io_addrout; // @[BuildingBlockNew.scala 296:22]
  assign ingress2_io_ctrl = instr3; // @[BuildingBlockNew.scala 165:20]
  assign middle_clock = clock;
  assign middle_io_in64_0 = ingress2_io_out64_0; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_1 = ingress2_io_out64_1; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_2 = ingress2_io_out64_2; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_3 = ingress2_io_out64_3; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_4 = ingress2_io_out64_4; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_5 = ingress2_io_out64_5; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_6 = ingress2_io_out64_6; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_7 = ingress2_io_out64_7; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_8 = ingress2_io_out64_8; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_9 = ingress2_io_out64_9; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_10 = ingress2_io_out64_10; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_11 = ingress2_io_out64_11; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_12 = ingress2_io_out64_12; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_13 = ingress2_io_out64_13; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_14 = ingress2_io_out64_14; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_15 = ingress2_io_out64_15; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_16 = ingress2_io_out64_16; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_17 = ingress2_io_out64_17; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_18 = ingress2_io_out64_18; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_19 = ingress2_io_out64_19; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_20 = ingress2_io_out64_20; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_21 = ingress2_io_out64_21; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_22 = ingress2_io_out64_22; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_23 = ingress2_io_out64_23; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_24 = ingress2_io_out64_24; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_25 = ingress2_io_out64_25; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_26 = ingress2_io_out64_26; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_27 = ingress2_io_out64_27; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_28 = ingress2_io_out64_28; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_29 = ingress2_io_out64_29; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_30 = ingress2_io_out64_30; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_31 = ingress2_io_out64_31; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_32 = ingress2_io_out64_32; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_33 = ingress2_io_out64_33; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_34 = ingress2_io_out64_34; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_35 = ingress2_io_out64_35; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_36 = ingress2_io_out64_36; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_37 = ingress2_io_out64_37; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_38 = ingress2_io_out64_38; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_39 = ingress2_io_out64_39; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_40 = ingress2_io_out64_40; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_41 = ingress2_io_out64_41; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_42 = ingress2_io_out64_42; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_43 = ingress2_io_out64_43; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_44 = ingress2_io_out64_44; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_45 = ingress2_io_out64_45; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_46 = ingress2_io_out64_46; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_47 = ingress2_io_out64_47; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_48 = ingress2_io_out64_48; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_49 = ingress2_io_out64_49; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_50 = ingress2_io_out64_50; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_51 = ingress2_io_out64_51; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_52 = ingress2_io_out64_52; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_53 = ingress2_io_out64_53; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_54 = ingress2_io_out64_54; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_55 = ingress2_io_out64_55; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_56 = ingress2_io_out64_56; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_57 = ingress2_io_out64_57; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_58 = ingress2_io_out64_58; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_59 = ingress2_io_out64_59; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_60 = ingress2_io_out64_60; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_61 = ingress2_io_out64_61; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_62 = ingress2_io_out64_62; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_63 = ingress2_io_out64_63; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_validin64_0 = ingress2_io_validout64_0; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_1 = ingress2_io_validout64_1; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_2 = ingress2_io_validout64_2; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_3 = ingress2_io_validout64_3; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_4 = ingress2_io_validout64_4; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_5 = ingress2_io_validout64_5; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_6 = ingress2_io_validout64_6; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_7 = ingress2_io_validout64_7; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_8 = ingress2_io_validout64_8; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_9 = ingress2_io_validout64_9; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_10 = ingress2_io_validout64_10; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_11 = ingress2_io_validout64_11; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_12 = ingress2_io_validout64_12; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_13 = ingress2_io_validout64_13; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_14 = ingress2_io_validout64_14; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_15 = ingress2_io_validout64_15; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_16 = ingress2_io_validout64_16; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_17 = ingress2_io_validout64_17; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_18 = ingress2_io_validout64_18; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_19 = ingress2_io_validout64_19; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_20 = ingress2_io_validout64_20; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_21 = ingress2_io_validout64_21; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_22 = ingress2_io_validout64_22; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_23 = ingress2_io_validout64_23; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_24 = ingress2_io_validout64_24; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_25 = ingress2_io_validout64_25; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_26 = ingress2_io_validout64_26; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_27 = ingress2_io_validout64_27; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_28 = ingress2_io_validout64_28; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_29 = ingress2_io_validout64_29; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_30 = ingress2_io_validout64_30; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_31 = ingress2_io_validout64_31; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_32 = ingress2_io_validout64_32; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_33 = ingress2_io_validout64_33; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_34 = ingress2_io_validout64_34; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_35 = ingress2_io_validout64_35; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_36 = ingress2_io_validout64_36; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_37 = ingress2_io_validout64_37; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_38 = ingress2_io_validout64_38; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_39 = ingress2_io_validout64_39; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_40 = ingress2_io_validout64_40; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_41 = ingress2_io_validout64_41; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_42 = ingress2_io_validout64_42; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_43 = ingress2_io_validout64_43; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_44 = ingress2_io_validout64_44; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_45 = ingress2_io_validout64_45; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_46 = ingress2_io_validout64_46; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_47 = ingress2_io_validout64_47; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_48 = ingress2_io_validout64_48; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_49 = ingress2_io_validout64_49; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_50 = ingress2_io_validout64_50; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_51 = ingress2_io_validout64_51; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_52 = ingress2_io_validout64_52; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_53 = ingress2_io_validout64_53; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_54 = ingress2_io_validout64_54; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_55 = ingress2_io_validout64_55; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_56 = ingress2_io_validout64_56; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_57 = ingress2_io_validout64_57; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_58 = ingress2_io_validout64_58; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_59 = ingress2_io_validout64_59; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_60 = ingress2_io_validout64_60; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_61 = ingress2_io_validout64_61; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_62 = ingress2_io_validout64_62; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_63 = ingress2_io_validout64_63; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_tagin_Tag = ingress2_io_tagout_Tag; // @[BuildingBlockNew.scala 299:19]
  assign middle_io_tagin_RoundCnt = ingress2_io_tagout_RoundCnt; // @[BuildingBlockNew.scala 299:19]
  assign middle_io_addrin = ingress2_io_addrout; // @[BuildingBlockNew.scala 300:20]
  assign middle_io_ctrl = instr4; // @[BuildingBlockNew.scala 166:18]
  assign egress1_clock = clock;
  assign egress1_io_in64_0 = middle_io_out64_0; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_1 = middle_io_out64_1; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_2 = middle_io_out64_2; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_3 = middle_io_out64_3; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_4 = middle_io_out64_4; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_5 = middle_io_out64_5; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_6 = middle_io_out64_6; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_7 = middle_io_out64_7; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_8 = middle_io_out64_8; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_9 = middle_io_out64_9; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_10 = middle_io_out64_10; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_11 = middle_io_out64_11; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_12 = middle_io_out64_12; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_13 = middle_io_out64_13; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_14 = middle_io_out64_14; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_15 = middle_io_out64_15; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_16 = middle_io_out64_16; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_17 = middle_io_out64_17; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_18 = middle_io_out64_18; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_19 = middle_io_out64_19; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_20 = middle_io_out64_20; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_21 = middle_io_out64_21; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_22 = middle_io_out64_22; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_23 = middle_io_out64_23; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_24 = middle_io_out64_24; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_25 = middle_io_out64_25; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_26 = middle_io_out64_26; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_27 = middle_io_out64_27; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_28 = middle_io_out64_28; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_29 = middle_io_out64_29; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_30 = middle_io_out64_30; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_31 = middle_io_out64_31; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_32 = middle_io_out64_32; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_33 = middle_io_out64_33; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_34 = middle_io_out64_34; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_35 = middle_io_out64_35; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_36 = middle_io_out64_36; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_37 = middle_io_out64_37; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_38 = middle_io_out64_38; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_39 = middle_io_out64_39; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_40 = middle_io_out64_40; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_41 = middle_io_out64_41; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_42 = middle_io_out64_42; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_43 = middle_io_out64_43; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_44 = middle_io_out64_44; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_45 = middle_io_out64_45; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_46 = middle_io_out64_46; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_47 = middle_io_out64_47; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_48 = middle_io_out64_48; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_49 = middle_io_out64_49; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_50 = middle_io_out64_50; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_51 = middle_io_out64_51; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_52 = middle_io_out64_52; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_53 = middle_io_out64_53; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_54 = middle_io_out64_54; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_55 = middle_io_out64_55; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_56 = middle_io_out64_56; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_57 = middle_io_out64_57; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_58 = middle_io_out64_58; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_59 = middle_io_out64_59; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_60 = middle_io_out64_60; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_61 = middle_io_out64_61; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_62 = middle_io_out64_62; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_63 = middle_io_out64_63; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_validin64_0 = middle_io_validout64_0; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_1 = middle_io_validout64_1; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_2 = middle_io_validout64_2; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_3 = middle_io_validout64_3; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_4 = middle_io_validout64_4; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_5 = middle_io_validout64_5; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_6 = middle_io_validout64_6; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_7 = middle_io_validout64_7; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_8 = middle_io_validout64_8; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_9 = middle_io_validout64_9; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_10 = middle_io_validout64_10; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_11 = middle_io_validout64_11; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_12 = middle_io_validout64_12; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_13 = middle_io_validout64_13; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_14 = middle_io_validout64_14; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_15 = middle_io_validout64_15; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_16 = middle_io_validout64_16; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_17 = middle_io_validout64_17; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_18 = middle_io_validout64_18; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_19 = middle_io_validout64_19; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_20 = middle_io_validout64_20; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_21 = middle_io_validout64_21; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_22 = middle_io_validout64_22; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_23 = middle_io_validout64_23; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_24 = middle_io_validout64_24; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_25 = middle_io_validout64_25; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_26 = middle_io_validout64_26; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_27 = middle_io_validout64_27; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_28 = middle_io_validout64_28; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_29 = middle_io_validout64_29; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_30 = middle_io_validout64_30; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_31 = middle_io_validout64_31; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_32 = middle_io_validout64_32; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_33 = middle_io_validout64_33; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_34 = middle_io_validout64_34; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_35 = middle_io_validout64_35; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_36 = middle_io_validout64_36; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_37 = middle_io_validout64_37; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_38 = middle_io_validout64_38; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_39 = middle_io_validout64_39; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_40 = middle_io_validout64_40; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_41 = middle_io_validout64_41; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_42 = middle_io_validout64_42; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_43 = middle_io_validout64_43; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_44 = middle_io_validout64_44; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_45 = middle_io_validout64_45; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_46 = middle_io_validout64_46; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_47 = middle_io_validout64_47; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_48 = middle_io_validout64_48; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_49 = middle_io_validout64_49; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_50 = middle_io_validout64_50; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_51 = middle_io_validout64_51; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_52 = middle_io_validout64_52; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_53 = middle_io_validout64_53; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_54 = middle_io_validout64_54; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_55 = middle_io_validout64_55; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_56 = middle_io_validout64_56; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_57 = middle_io_validout64_57; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_58 = middle_io_validout64_58; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_59 = middle_io_validout64_59; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_60 = middle_io_validout64_60; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_61 = middle_io_validout64_61; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_62 = middle_io_validout64_62; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_63 = middle_io_validout64_63; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_tagin_Tag = middle_io_tagout_Tag; // @[BuildingBlockNew.scala 303:20]
  assign egress1_io_tagin_RoundCnt = middle_io_tagout_RoundCnt; // @[BuildingBlockNew.scala 303:20]
  assign egress1_io_addrin = middle_io_addrout; // @[BuildingBlockNew.scala 304:21]
  assign egress1_io_ctrl = instr5; // @[BuildingBlockNew.scala 167:19]
  assign egress2_clock = clock;
  assign egress2_io_in64_0 = egress1_io_out64_0; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_1 = egress1_io_out64_1; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_2 = egress1_io_out64_2; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_3 = egress1_io_out64_3; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_4 = egress1_io_out64_4; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_5 = egress1_io_out64_5; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_6 = egress1_io_out64_6; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_7 = egress1_io_out64_7; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_8 = egress1_io_out64_8; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_9 = egress1_io_out64_9; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_10 = egress1_io_out64_10; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_11 = egress1_io_out64_11; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_12 = egress1_io_out64_12; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_13 = egress1_io_out64_13; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_14 = egress1_io_out64_14; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_15 = egress1_io_out64_15; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_16 = egress1_io_out64_16; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_17 = egress1_io_out64_17; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_18 = egress1_io_out64_18; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_19 = egress1_io_out64_19; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_20 = egress1_io_out64_20; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_21 = egress1_io_out64_21; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_22 = egress1_io_out64_22; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_23 = egress1_io_out64_23; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_24 = egress1_io_out64_24; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_25 = egress1_io_out64_25; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_26 = egress1_io_out64_26; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_27 = egress1_io_out64_27; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_28 = egress1_io_out64_28; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_29 = egress1_io_out64_29; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_30 = egress1_io_out64_30; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_31 = egress1_io_out64_31; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_32 = egress1_io_out64_32; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_33 = egress1_io_out64_33; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_34 = egress1_io_out64_34; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_35 = egress1_io_out64_35; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_36 = egress1_io_out64_36; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_37 = egress1_io_out64_37; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_38 = egress1_io_out64_38; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_39 = egress1_io_out64_39; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_40 = egress1_io_out64_40; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_41 = egress1_io_out64_41; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_42 = egress1_io_out64_42; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_43 = egress1_io_out64_43; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_44 = egress1_io_out64_44; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_45 = egress1_io_out64_45; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_46 = egress1_io_out64_46; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_47 = egress1_io_out64_47; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_48 = egress1_io_out64_48; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_49 = egress1_io_out64_49; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_50 = egress1_io_out64_50; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_51 = egress1_io_out64_51; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_52 = egress1_io_out64_52; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_53 = egress1_io_out64_53; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_54 = egress1_io_out64_54; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_55 = egress1_io_out64_55; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_56 = egress1_io_out64_56; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_57 = egress1_io_out64_57; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_58 = egress1_io_out64_58; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_59 = egress1_io_out64_59; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_60 = egress1_io_out64_60; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_61 = egress1_io_out64_61; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_62 = egress1_io_out64_62; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_63 = egress1_io_out64_63; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_validin64_0 = egress1_io_validout64_0; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_1 = egress1_io_validout64_1; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_2 = egress1_io_validout64_2; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_3 = egress1_io_validout64_3; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_4 = egress1_io_validout64_4; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_5 = egress1_io_validout64_5; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_6 = egress1_io_validout64_6; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_7 = egress1_io_validout64_7; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_8 = egress1_io_validout64_8; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_9 = egress1_io_validout64_9; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_10 = egress1_io_validout64_10; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_11 = egress1_io_validout64_11; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_12 = egress1_io_validout64_12; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_13 = egress1_io_validout64_13; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_14 = egress1_io_validout64_14; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_15 = egress1_io_validout64_15; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_16 = egress1_io_validout64_16; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_17 = egress1_io_validout64_17; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_18 = egress1_io_validout64_18; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_19 = egress1_io_validout64_19; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_20 = egress1_io_validout64_20; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_21 = egress1_io_validout64_21; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_22 = egress1_io_validout64_22; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_23 = egress1_io_validout64_23; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_24 = egress1_io_validout64_24; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_25 = egress1_io_validout64_25; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_26 = egress1_io_validout64_26; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_27 = egress1_io_validout64_27; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_28 = egress1_io_validout64_28; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_29 = egress1_io_validout64_29; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_30 = egress1_io_validout64_30; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_31 = egress1_io_validout64_31; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_32 = egress1_io_validout64_32; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_33 = egress1_io_validout64_33; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_34 = egress1_io_validout64_34; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_35 = egress1_io_validout64_35; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_36 = egress1_io_validout64_36; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_37 = egress1_io_validout64_37; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_38 = egress1_io_validout64_38; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_39 = egress1_io_validout64_39; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_40 = egress1_io_validout64_40; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_41 = egress1_io_validout64_41; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_42 = egress1_io_validout64_42; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_43 = egress1_io_validout64_43; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_44 = egress1_io_validout64_44; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_45 = egress1_io_validout64_45; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_46 = egress1_io_validout64_46; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_47 = egress1_io_validout64_47; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_48 = egress1_io_validout64_48; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_49 = egress1_io_validout64_49; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_50 = egress1_io_validout64_50; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_51 = egress1_io_validout64_51; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_52 = egress1_io_validout64_52; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_53 = egress1_io_validout64_53; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_54 = egress1_io_validout64_54; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_55 = egress1_io_validout64_55; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_56 = egress1_io_validout64_56; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_57 = egress1_io_validout64_57; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_58 = egress1_io_validout64_58; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_59 = egress1_io_validout64_59; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_60 = egress1_io_validout64_60; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_61 = egress1_io_validout64_61; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_62 = egress1_io_validout64_62; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_63 = egress1_io_validout64_63; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_tagin_Tag = egress1_io_tagout_Tag; // @[BuildingBlockNew.scala 307:20]
  assign egress2_io_tagin_RoundCnt = egress1_io_tagout_RoundCnt; // @[BuildingBlockNew.scala 307:20]
  assign egress2_io_addrin = egress1_io_addrout; // @[BuildingBlockNew.scala 308:21]
  assign egress2_io_ctrl = instr6; // @[BuildingBlockNew.scala 168:19]
  always @(posedge clock) begin
    if (reset) begin // @[BuildingBlockNew.scala 40:20]
      PC1 <= 8'h0; // @[BuildingBlockNew.scala 40:20]
    end else begin
      PC1 <= io_PC1_in; // @[BuildingBlockNew.scala 154:7]
    end
    if (reset) begin // @[BuildingBlockNew.scala 41:20]
      PC2 <= 8'h0; // @[BuildingBlockNew.scala 41:20]
    end else begin
      PC2 <= PC1; // @[BuildingBlockNew.scala 155:7]
    end
    if (reset) begin // @[BuildingBlockNew.scala 42:20]
      PC3 <= 8'h0; // @[BuildingBlockNew.scala 42:20]
    end else begin
      PC3 <= PC2; // @[BuildingBlockNew.scala 156:7]
    end
    if (reset) begin // @[BuildingBlockNew.scala 43:20]
      PC4 <= 8'h0; // @[BuildingBlockNew.scala 43:20]
    end else begin
      PC4 <= PC3; // @[BuildingBlockNew.scala 157:7]
    end
    if (reset) begin // @[BuildingBlockNew.scala 44:20]
      PC5 <= 8'h0; // @[BuildingBlockNew.scala 44:20]
    end else begin
      PC5 <= PC4; // @[BuildingBlockNew.scala 158:7]
    end
    if (reset) begin // @[BuildingBlockNew.scala 45:20]
      PC6 <= 8'h0; // @[BuildingBlockNew.scala 45:20]
    end else begin
      PC6 <= PC5; // @[BuildingBlockNew.scala 159:7]
    end
    if (reset) begin // @[BuildingBlockNew.scala 46:24]
      wrAddr1 <= 8'h0; // @[BuildingBlockNew.scala 46:24]
    end else if (io_wr_en_mem1) begin // @[BuildingBlockNew.scala 223:22]
      wrAddr1 <= _wrAddr1_T_1; // @[BuildingBlockNew.scala 226:13]
    end
    if (reset) begin // @[BuildingBlockNew.scala 47:24]
      wrAddr2 <= 8'h0; // @[BuildingBlockNew.scala 47:24]
    end else if (io_wr_en_mem2) begin // @[BuildingBlockNew.scala 232:22]
      wrAddr2 <= _wrAddr2_T_1; // @[BuildingBlockNew.scala 235:13]
    end
    if (reset) begin // @[BuildingBlockNew.scala 48:24]
      wrAddr3 <= 8'h0; // @[BuildingBlockNew.scala 48:24]
    end else if (io_wr_en_mem3) begin // @[BuildingBlockNew.scala 241:22]
      wrAddr3 <= _wrAddr3_T_1; // @[BuildingBlockNew.scala 244:13]
    end
    if (reset) begin // @[BuildingBlockNew.scala 49:24]
      wrAddr4 <= 8'h0; // @[BuildingBlockNew.scala 49:24]
    end else if (io_wr_en_mem4) begin // @[BuildingBlockNew.scala 250:22]
      wrAddr4 <= _wrAddr4_T_1; // @[BuildingBlockNew.scala 253:13]
    end
    if (reset) begin // @[BuildingBlockNew.scala 50:24]
      wrAddr5 <= 8'h0; // @[BuildingBlockNew.scala 50:24]
    end else if (io_wr_en_mem5) begin // @[BuildingBlockNew.scala 259:22]
      wrAddr5 <= _wrAddr5_T_1; // @[BuildingBlockNew.scala 262:13]
    end
    if (reset) begin // @[BuildingBlockNew.scala 51:24]
      wrAddr6 <= 8'h0; // @[BuildingBlockNew.scala 51:24]
    end else if (io_wr_en_mem6) begin // @[BuildingBlockNew.scala 268:22]
      wrAddr6 <= _wrAddr6_T_1; // @[BuildingBlockNew.scala 271:13]
    end
    instr1 <= Mem1_R0_data; // @[BuildingBlockNew.scala 223:22 BuildingBlockNew.scala 229:12]
    instr2 <= Mem2_R0_data; // @[BuildingBlockNew.scala 232:22 BuildingBlockNew.scala 238:12]
    instr3 <= Mem3_R0_data; // @[BuildingBlockNew.scala 241:22 BuildingBlockNew.scala 247:12]
    instr4 <= Mem4_R0_data; // @[BuildingBlockNew.scala 250:22 BuildingBlockNew.scala 256:12]
    instr5 <= Mem5_R0_data; // @[BuildingBlockNew.scala 259:22 BuildingBlockNew.scala 265:12]
    instr6 <= Mem6_R0_data; // @[BuildingBlockNew.scala 268:22 BuildingBlockNew.scala 274:12]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  PC1 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  PC2 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  PC3 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  PC4 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  PC5 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  PC6 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  wrAddr1 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  wrAddr2 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  wrAddr3 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  wrAddr4 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  wrAddr5 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  wrAddr6 = _RAND_11[7:0];
  _RAND_12 = {9{`RANDOM}};
  instr1 = _RAND_12[287:0];
  _RAND_13 = {4{`RANDOM}};
  instr2 = _RAND_13[127:0];
  _RAND_14 = {4{`RANDOM}};
  instr3 = _RAND_14[127:0];
  _RAND_15 = {4{`RANDOM}};
  instr4 = _RAND_15[127:0];
  _RAND_16 = {4{`RANDOM}};
  instr5 = _RAND_16[127:0];
  _RAND_17 = {4{`RANDOM}};
  instr6 = _RAND_17[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PEArray(
  input          clock,
  input          reset,
  input          io_wr_en_mem1_0,
  input          io_wr_en_mem1_1,
  input          io_wr_en_mem1_2,
  input          io_wr_en_mem1_3,
  input          io_wr_en_mem1_4,
  input          io_wr_en_mem1_5,
  input          io_wr_en_mem1_6,
  input          io_wr_en_mem1_7,
  input          io_wr_en_mem1_8,
  input          io_wr_en_mem1_9,
  input          io_wr_en_mem1_10,
  input          io_wr_en_mem1_11,
  input          io_wr_en_mem1_12,
  input          io_wr_en_mem1_13,
  input          io_wr_en_mem1_14,
  input          io_wr_en_mem1_15,
  input          io_wr_en_mem2_0,
  input          io_wr_en_mem2_1,
  input          io_wr_en_mem2_2,
  input          io_wr_en_mem2_3,
  input          io_wr_en_mem2_4,
  input          io_wr_en_mem2_5,
  input          io_wr_en_mem2_6,
  input          io_wr_en_mem2_7,
  input          io_wr_en_mem2_8,
  input          io_wr_en_mem2_9,
  input          io_wr_en_mem2_10,
  input          io_wr_en_mem2_11,
  input          io_wr_en_mem2_12,
  input          io_wr_en_mem2_13,
  input          io_wr_en_mem2_14,
  input          io_wr_en_mem2_15,
  input          io_wr_en_mem3_0,
  input          io_wr_en_mem3_1,
  input          io_wr_en_mem3_2,
  input          io_wr_en_mem3_3,
  input          io_wr_en_mem3_4,
  input          io_wr_en_mem3_5,
  input          io_wr_en_mem3_6,
  input          io_wr_en_mem3_7,
  input          io_wr_en_mem3_8,
  input          io_wr_en_mem3_9,
  input          io_wr_en_mem3_10,
  input          io_wr_en_mem3_11,
  input          io_wr_en_mem3_12,
  input          io_wr_en_mem3_13,
  input          io_wr_en_mem3_14,
  input          io_wr_en_mem3_15,
  input          io_wr_en_mem4_0,
  input          io_wr_en_mem4_1,
  input          io_wr_en_mem4_2,
  input          io_wr_en_mem4_3,
  input          io_wr_en_mem4_4,
  input          io_wr_en_mem4_5,
  input          io_wr_en_mem4_6,
  input          io_wr_en_mem4_7,
  input          io_wr_en_mem4_8,
  input          io_wr_en_mem4_9,
  input          io_wr_en_mem4_10,
  input          io_wr_en_mem4_11,
  input          io_wr_en_mem4_12,
  input          io_wr_en_mem4_13,
  input          io_wr_en_mem4_14,
  input          io_wr_en_mem4_15,
  input          io_wr_en_mem5_0,
  input          io_wr_en_mem5_1,
  input          io_wr_en_mem5_2,
  input          io_wr_en_mem5_3,
  input          io_wr_en_mem5_4,
  input          io_wr_en_mem5_5,
  input          io_wr_en_mem5_6,
  input          io_wr_en_mem5_7,
  input          io_wr_en_mem5_8,
  input          io_wr_en_mem5_9,
  input          io_wr_en_mem5_10,
  input          io_wr_en_mem5_11,
  input          io_wr_en_mem5_12,
  input          io_wr_en_mem5_13,
  input          io_wr_en_mem5_14,
  input          io_wr_en_mem5_15,
  input          io_wr_en_mem6_0,
  input          io_wr_en_mem6_1,
  input          io_wr_en_mem6_2,
  input          io_wr_en_mem6_3,
  input          io_wr_en_mem6_4,
  input          io_wr_en_mem6_5,
  input          io_wr_en_mem6_6,
  input          io_wr_en_mem6_7,
  input          io_wr_en_mem6_8,
  input          io_wr_en_mem6_9,
  input          io_wr_en_mem6_10,
  input          io_wr_en_mem6_11,
  input          io_wr_en_mem6_12,
  input          io_wr_en_mem6_13,
  input          io_wr_en_mem6_14,
  input          io_wr_en_mem6_15,
  input  [287:0] io_wr_instr_mem1_0,
  input  [287:0] io_wr_instr_mem1_1,
  input  [287:0] io_wr_instr_mem1_2,
  input  [287:0] io_wr_instr_mem1_3,
  input  [287:0] io_wr_instr_mem1_4,
  input  [287:0] io_wr_instr_mem1_5,
  input  [287:0] io_wr_instr_mem1_6,
  input  [287:0] io_wr_instr_mem1_7,
  input  [287:0] io_wr_instr_mem1_8,
  input  [287:0] io_wr_instr_mem1_9,
  input  [287:0] io_wr_instr_mem1_10,
  input  [287:0] io_wr_instr_mem1_11,
  input  [287:0] io_wr_instr_mem1_12,
  input  [287:0] io_wr_instr_mem1_13,
  input  [287:0] io_wr_instr_mem1_14,
  input  [287:0] io_wr_instr_mem1_15,
  input  [127:0] io_wr_instr_mem2_0,
  input  [127:0] io_wr_instr_mem2_1,
  input  [127:0] io_wr_instr_mem2_2,
  input  [127:0] io_wr_instr_mem2_3,
  input  [127:0] io_wr_instr_mem2_4,
  input  [127:0] io_wr_instr_mem2_5,
  input  [127:0] io_wr_instr_mem2_6,
  input  [127:0] io_wr_instr_mem2_7,
  input  [127:0] io_wr_instr_mem2_8,
  input  [127:0] io_wr_instr_mem2_9,
  input  [127:0] io_wr_instr_mem2_10,
  input  [127:0] io_wr_instr_mem2_11,
  input  [127:0] io_wr_instr_mem2_12,
  input  [127:0] io_wr_instr_mem2_13,
  input  [127:0] io_wr_instr_mem2_14,
  input  [127:0] io_wr_instr_mem2_15,
  input  [127:0] io_wr_instr_mem3_0,
  input  [127:0] io_wr_instr_mem3_1,
  input  [127:0] io_wr_instr_mem3_2,
  input  [127:0] io_wr_instr_mem3_3,
  input  [127:0] io_wr_instr_mem3_4,
  input  [127:0] io_wr_instr_mem3_5,
  input  [127:0] io_wr_instr_mem3_6,
  input  [127:0] io_wr_instr_mem3_7,
  input  [127:0] io_wr_instr_mem3_8,
  input  [127:0] io_wr_instr_mem3_9,
  input  [127:0] io_wr_instr_mem3_10,
  input  [127:0] io_wr_instr_mem3_11,
  input  [127:0] io_wr_instr_mem3_12,
  input  [127:0] io_wr_instr_mem3_13,
  input  [127:0] io_wr_instr_mem3_14,
  input  [127:0] io_wr_instr_mem3_15,
  input  [127:0] io_wr_instr_mem4_0,
  input  [127:0] io_wr_instr_mem4_1,
  input  [127:0] io_wr_instr_mem4_2,
  input  [127:0] io_wr_instr_mem4_3,
  input  [127:0] io_wr_instr_mem4_4,
  input  [127:0] io_wr_instr_mem4_5,
  input  [127:0] io_wr_instr_mem4_6,
  input  [127:0] io_wr_instr_mem4_7,
  input  [127:0] io_wr_instr_mem4_8,
  input  [127:0] io_wr_instr_mem4_9,
  input  [127:0] io_wr_instr_mem4_10,
  input  [127:0] io_wr_instr_mem4_11,
  input  [127:0] io_wr_instr_mem4_12,
  input  [127:0] io_wr_instr_mem4_13,
  input  [127:0] io_wr_instr_mem4_14,
  input  [127:0] io_wr_instr_mem4_15,
  input  [127:0] io_wr_instr_mem5_0,
  input  [127:0] io_wr_instr_mem5_1,
  input  [127:0] io_wr_instr_mem5_2,
  input  [127:0] io_wr_instr_mem5_3,
  input  [127:0] io_wr_instr_mem5_4,
  input  [127:0] io_wr_instr_mem5_5,
  input  [127:0] io_wr_instr_mem5_6,
  input  [127:0] io_wr_instr_mem5_7,
  input  [127:0] io_wr_instr_mem5_8,
  input  [127:0] io_wr_instr_mem5_9,
  input  [127:0] io_wr_instr_mem5_10,
  input  [127:0] io_wr_instr_mem5_11,
  input  [127:0] io_wr_instr_mem5_12,
  input  [127:0] io_wr_instr_mem5_13,
  input  [127:0] io_wr_instr_mem5_14,
  input  [127:0] io_wr_instr_mem5_15,
  input  [127:0] io_wr_instr_mem6_0,
  input  [127:0] io_wr_instr_mem6_1,
  input  [127:0] io_wr_instr_mem6_2,
  input  [127:0] io_wr_instr_mem6_3,
  input  [127:0] io_wr_instr_mem6_4,
  input  [127:0] io_wr_instr_mem6_5,
  input  [127:0] io_wr_instr_mem6_6,
  input  [127:0] io_wr_instr_mem6_7,
  input  [127:0] io_wr_instr_mem6_8,
  input  [127:0] io_wr_instr_mem6_9,
  input  [127:0] io_wr_instr_mem6_10,
  input  [127:0] io_wr_instr_mem6_11,
  input  [127:0] io_wr_instr_mem6_12,
  input  [127:0] io_wr_instr_mem6_13,
  input  [127:0] io_wr_instr_mem6_14,
  input  [127:0] io_wr_instr_mem6_15,
  input  [63:0]  io_d_in_0_a,
  input          io_d_in_0_valid_a,
  input  [63:0]  io_d_in_0_b,
  input          io_d_in_0_valid_b,
  input  [63:0]  io_d_in_1_a,
  input          io_d_in_1_valid_a,
  input  [63:0]  io_d_in_1_b,
  input          io_d_in_1_valid_b,
  input  [63:0]  io_d_in_2_a,
  input          io_d_in_2_valid_a,
  input  [63:0]  io_d_in_2_b,
  input          io_d_in_2_valid_b,
  input  [63:0]  io_d_in_3_a,
  input          io_d_in_3_valid_a,
  input  [63:0]  io_d_in_3_b,
  input          io_d_in_3_valid_b,
  input  [63:0]  io_d_in_4_a,
  input          io_d_in_4_valid_a,
  input  [63:0]  io_d_in_4_b,
  input          io_d_in_4_valid_b,
  input  [63:0]  io_d_in_5_a,
  input          io_d_in_5_valid_a,
  input  [63:0]  io_d_in_5_b,
  input          io_d_in_5_valid_b,
  input  [63:0]  io_d_in_6_a,
  input          io_d_in_6_valid_a,
  input  [63:0]  io_d_in_6_b,
  input          io_d_in_6_valid_b,
  input  [63:0]  io_d_in_7_a,
  input          io_d_in_7_valid_a,
  input  [63:0]  io_d_in_7_b,
  input          io_d_in_7_valid_b,
  input  [63:0]  io_d_in_8_a,
  input          io_d_in_8_valid_a,
  input  [63:0]  io_d_in_8_b,
  input          io_d_in_8_valid_b,
  input  [63:0]  io_d_in_9_a,
  input          io_d_in_9_valid_a,
  input  [63:0]  io_d_in_9_b,
  input          io_d_in_9_valid_b,
  input  [63:0]  io_d_in_10_a,
  input          io_d_in_10_valid_a,
  input  [63:0]  io_d_in_10_b,
  input          io_d_in_10_valid_b,
  input  [63:0]  io_d_in_11_a,
  input          io_d_in_11_valid_a,
  input  [63:0]  io_d_in_11_b,
  input          io_d_in_11_valid_b,
  input  [63:0]  io_d_in_12_a,
  input          io_d_in_12_valid_a,
  input  [63:0]  io_d_in_12_b,
  input          io_d_in_12_valid_b,
  input  [63:0]  io_d_in_13_a,
  input          io_d_in_13_valid_a,
  input  [63:0]  io_d_in_13_b,
  input          io_d_in_13_valid_b,
  input  [63:0]  io_d_in_14_a,
  input          io_d_in_14_valid_a,
  input  [63:0]  io_d_in_14_b,
  input          io_d_in_14_valid_b,
  input  [63:0]  io_d_in_15_a,
  input          io_d_in_15_valid_a,
  input  [63:0]  io_d_in_15_b,
  input          io_d_in_15_valid_b,
  input  [63:0]  io_d_in_16_a,
  input          io_d_in_16_valid_a,
  input  [63:0]  io_d_in_16_b,
  input          io_d_in_16_valid_b,
  input  [63:0]  io_d_in_17_a,
  input          io_d_in_17_valid_a,
  input  [63:0]  io_d_in_17_b,
  input          io_d_in_17_valid_b,
  input  [63:0]  io_d_in_18_a,
  input          io_d_in_18_valid_a,
  input  [63:0]  io_d_in_18_b,
  input          io_d_in_18_valid_b,
  input  [63:0]  io_d_in_19_a,
  input          io_d_in_19_valid_a,
  input  [63:0]  io_d_in_19_b,
  input          io_d_in_19_valid_b,
  input  [63:0]  io_d_in_20_a,
  input          io_d_in_20_valid_a,
  input  [63:0]  io_d_in_20_b,
  input          io_d_in_20_valid_b,
  input  [63:0]  io_d_in_21_a,
  input          io_d_in_21_valid_a,
  input  [63:0]  io_d_in_21_b,
  input          io_d_in_21_valid_b,
  input  [63:0]  io_d_in_22_a,
  input          io_d_in_22_valid_a,
  input  [63:0]  io_d_in_22_b,
  input          io_d_in_22_valid_b,
  input  [63:0]  io_d_in_23_a,
  input          io_d_in_23_valid_a,
  input  [63:0]  io_d_in_23_b,
  input          io_d_in_23_valid_b,
  input  [63:0]  io_d_in_24_a,
  input          io_d_in_24_valid_a,
  input  [63:0]  io_d_in_24_b,
  input          io_d_in_24_valid_b,
  input  [63:0]  io_d_in_25_a,
  input          io_d_in_25_valid_a,
  input  [63:0]  io_d_in_25_b,
  input          io_d_in_25_valid_b,
  input  [63:0]  io_d_in_26_a,
  input          io_d_in_26_valid_a,
  input  [63:0]  io_d_in_26_b,
  input          io_d_in_26_valid_b,
  input  [63:0]  io_d_in_27_a,
  input          io_d_in_27_valid_a,
  input  [63:0]  io_d_in_27_b,
  input          io_d_in_27_valid_b,
  input  [63:0]  io_d_in_28_a,
  input          io_d_in_28_valid_a,
  input  [63:0]  io_d_in_28_b,
  input          io_d_in_28_valid_b,
  input  [63:0]  io_d_in_29_a,
  input          io_d_in_29_valid_a,
  input  [63:0]  io_d_in_29_b,
  input          io_d_in_29_valid_b,
  input  [63:0]  io_d_in_30_a,
  input          io_d_in_30_valid_a,
  input  [63:0]  io_d_in_30_b,
  input          io_d_in_30_valid_b,
  input  [63:0]  io_d_in_31_a,
  input          io_d_in_31_valid_a,
  input  [63:0]  io_d_in_31_b,
  input          io_d_in_31_valid_b,
  output [63:0]  io_d_out_0_a,
  output         io_d_out_0_valid_a,
  output [63:0]  io_d_out_0_b,
  output         io_d_out_0_valid_b,
  output [63:0]  io_d_out_1_a,
  output         io_d_out_1_valid_a,
  output [63:0]  io_d_out_1_b,
  output         io_d_out_1_valid_b,
  output [63:0]  io_d_out_2_a,
  output         io_d_out_2_valid_a,
  output [63:0]  io_d_out_2_b,
  output         io_d_out_2_valid_b,
  output [63:0]  io_d_out_3_a,
  output         io_d_out_3_valid_a,
  output [63:0]  io_d_out_3_b,
  output         io_d_out_3_valid_b,
  output [63:0]  io_d_out_4_a,
  output         io_d_out_4_valid_a,
  output [63:0]  io_d_out_4_b,
  output         io_d_out_4_valid_b,
  output [63:0]  io_d_out_5_a,
  output         io_d_out_5_valid_a,
  output [63:0]  io_d_out_5_b,
  output         io_d_out_5_valid_b,
  output [63:0]  io_d_out_6_a,
  output         io_d_out_6_valid_a,
  output [63:0]  io_d_out_6_b,
  output         io_d_out_6_valid_b,
  output [63:0]  io_d_out_7_a,
  output         io_d_out_7_valid_a,
  output [63:0]  io_d_out_7_b,
  output         io_d_out_7_valid_b,
  output [63:0]  io_d_out_8_a,
  output         io_d_out_8_valid_a,
  output [63:0]  io_d_out_8_b,
  output         io_d_out_8_valid_b,
  output [63:0]  io_d_out_9_a,
  output         io_d_out_9_valid_a,
  output [63:0]  io_d_out_9_b,
  output         io_d_out_9_valid_b,
  output [63:0]  io_d_out_10_a,
  output         io_d_out_10_valid_a,
  output [63:0]  io_d_out_10_b,
  output         io_d_out_10_valid_b,
  output [63:0]  io_d_out_11_a,
  output         io_d_out_11_valid_a,
  output [63:0]  io_d_out_11_b,
  output         io_d_out_11_valid_b,
  output [63:0]  io_d_out_12_a,
  output         io_d_out_12_valid_a,
  output [63:0]  io_d_out_12_b,
  output         io_d_out_12_valid_b,
  output [63:0]  io_d_out_13_a,
  output         io_d_out_13_valid_a,
  output [63:0]  io_d_out_13_b,
  output         io_d_out_13_valid_b,
  output [63:0]  io_d_out_14_a,
  output         io_d_out_14_valid_a,
  output [63:0]  io_d_out_14_b,
  output         io_d_out_14_valid_b,
  output [63:0]  io_d_out_15_a,
  output         io_d_out_15_valid_a,
  output [63:0]  io_d_out_15_b,
  output         io_d_out_15_valid_b,
  output [63:0]  io_d_out_16_a,
  output         io_d_out_16_valid_a,
  output [63:0]  io_d_out_16_b,
  output         io_d_out_16_valid_b,
  output [63:0]  io_d_out_17_a,
  output         io_d_out_17_valid_a,
  output [63:0]  io_d_out_17_b,
  output         io_d_out_17_valid_b,
  output [63:0]  io_d_out_18_a,
  output         io_d_out_18_valid_a,
  output [63:0]  io_d_out_18_b,
  output         io_d_out_18_valid_b,
  output [63:0]  io_d_out_19_a,
  output         io_d_out_19_valid_a,
  output [63:0]  io_d_out_19_b,
  output         io_d_out_19_valid_b,
  output [63:0]  io_d_out_20_a,
  output         io_d_out_20_valid_a,
  output [63:0]  io_d_out_20_b,
  output         io_d_out_20_valid_b,
  output [63:0]  io_d_out_21_a,
  output         io_d_out_21_valid_a,
  output [63:0]  io_d_out_21_b,
  output         io_d_out_21_valid_b,
  output [63:0]  io_d_out_22_a,
  output         io_d_out_22_valid_a,
  output [63:0]  io_d_out_22_b,
  output         io_d_out_22_valid_b,
  output [63:0]  io_d_out_23_a,
  output         io_d_out_23_valid_a,
  output [63:0]  io_d_out_23_b,
  output         io_d_out_23_valid_b,
  output [63:0]  io_d_out_24_a,
  output         io_d_out_24_valid_a,
  output [63:0]  io_d_out_24_b,
  output         io_d_out_24_valid_b,
  output [63:0]  io_d_out_25_a,
  output         io_d_out_25_valid_a,
  output [63:0]  io_d_out_25_b,
  output         io_d_out_25_valid_b,
  output [63:0]  io_d_out_26_a,
  output         io_d_out_26_valid_a,
  output [63:0]  io_d_out_26_b,
  output         io_d_out_26_valid_b,
  output [63:0]  io_d_out_27_a,
  output         io_d_out_27_valid_a,
  output [63:0]  io_d_out_27_b,
  output         io_d_out_27_valid_b,
  output [63:0]  io_d_out_28_a,
  output         io_d_out_28_valid_a,
  output [63:0]  io_d_out_28_b,
  output         io_d_out_28_valid_b,
  output [63:0]  io_d_out_29_a,
  output         io_d_out_29_valid_a,
  output [63:0]  io_d_out_29_b,
  output         io_d_out_29_valid_b,
  output [63:0]  io_d_out_30_a,
  output         io_d_out_30_valid_a,
  output [63:0]  io_d_out_30_b,
  output         io_d_out_30_valid_b,
  output [63:0]  io_d_out_31_a,
  output         io_d_out_31_valid_a,
  output [63:0]  io_d_out_31_b,
  output         io_d_out_31_valid_b,
  input  [1:0]   io_Tag_in_Tag,
  input  [2:0]   io_Tag_in_RoundCnt,
  output [1:0]   io_Tag_out_Tag,
  output [2:0]   io_Tag_out_RoundCnt,
  input  [7:0]   io_Addr_in,
  output [7:0]   io_Addr_out,
  input  [7:0]   io_PC_in,
  output [7:0]   io_PC_out,
  input          io_beginRun
);
  wire  array_0_clock; // @[Array.scala 41:54]
  wire  array_0_reset; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_0_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_0_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_0_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_0_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_0_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_0_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_0_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_0_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_0_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_0_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_0_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_0_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_0_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_0_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_0_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_0_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_0_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_0_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_0_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_0_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_0_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_0_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_0_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_0_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_1_clock; // @[Array.scala 41:54]
  wire  array_1_reset; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_1_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_1_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_1_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_1_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_1_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_1_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_1_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_1_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_1_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_1_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_1_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_1_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_1_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_1_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_1_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_1_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_1_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_1_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_1_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_1_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_1_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_1_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_1_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_1_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_2_clock; // @[Array.scala 41:54]
  wire  array_2_reset; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_2_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_2_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_2_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_2_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_2_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_2_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_2_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_2_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_2_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_2_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_2_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_2_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_2_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_2_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_2_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_2_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_2_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_2_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_2_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_2_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_2_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_2_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_2_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_2_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_3_clock; // @[Array.scala 41:54]
  wire  array_3_reset; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_3_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_3_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_3_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_3_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_3_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_3_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_3_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_3_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_3_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_3_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_3_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_3_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_3_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_3_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_3_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_3_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_3_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_3_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_3_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_3_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_3_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_3_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_3_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_3_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_4_clock; // @[Array.scala 41:54]
  wire  array_4_reset; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_4_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_4_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_4_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_4_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_4_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_4_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_4_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_4_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_4_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_4_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_4_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_4_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_4_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_4_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_4_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_4_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_4_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_4_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_4_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_4_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_4_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_4_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_4_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_4_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_5_clock; // @[Array.scala 41:54]
  wire  array_5_reset; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_5_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_5_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_5_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_5_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_5_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_5_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_5_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_5_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_5_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_5_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_5_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_5_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_5_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_5_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_5_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_5_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_5_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_5_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_5_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_5_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_5_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_5_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_5_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_5_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_6_clock; // @[Array.scala 41:54]
  wire  array_6_reset; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_6_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_6_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_6_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_6_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_6_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_6_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_6_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_6_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_6_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_6_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_6_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_6_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_6_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_6_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_6_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_6_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_6_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_6_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_6_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_6_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_6_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_6_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_6_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_6_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_7_clock; // @[Array.scala 41:54]
  wire  array_7_reset; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_7_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_7_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_7_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_7_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_7_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_7_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_7_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_7_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_7_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_7_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_7_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_7_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_7_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_7_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_7_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_7_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_7_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_7_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_7_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_7_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_7_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_7_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_7_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_7_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_8_clock; // @[Array.scala 41:54]
  wire  array_8_reset; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_8_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_8_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_8_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_8_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_8_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_8_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_8_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_8_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_8_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_8_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_8_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_8_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_8_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_8_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_8_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_8_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_8_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_8_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_8_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_8_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_8_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_8_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_8_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_8_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_9_clock; // @[Array.scala 41:54]
  wire  array_9_reset; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_9_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_9_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_9_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_9_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_9_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_9_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_9_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_9_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_9_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_9_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_9_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_9_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_9_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_9_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_9_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_9_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_9_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_9_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_9_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_9_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_9_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_9_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_9_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_9_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_10_clock; // @[Array.scala 41:54]
  wire  array_10_reset; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_10_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_10_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_10_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_10_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_10_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_10_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_10_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_10_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_10_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_10_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_10_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_10_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_10_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_10_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_10_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_10_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_10_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_10_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_10_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_10_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_10_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_10_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_10_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_10_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_11_clock; // @[Array.scala 41:54]
  wire  array_11_reset; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_11_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_11_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_11_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_11_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_11_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_11_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_11_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_11_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_11_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_11_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_11_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_11_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_11_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_11_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_11_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_11_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_11_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_11_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_11_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_11_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_11_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_11_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_11_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_11_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_12_clock; // @[Array.scala 41:54]
  wire  array_12_reset; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_12_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_12_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_12_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_12_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_12_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_12_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_12_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_12_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_12_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_12_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_12_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_12_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_12_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_12_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_12_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_12_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_12_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_12_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_12_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_12_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_12_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_12_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_12_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_12_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_13_clock; // @[Array.scala 41:54]
  wire  array_13_reset; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_13_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_13_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_13_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_13_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_13_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_13_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_13_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_13_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_13_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_13_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_13_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_13_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_13_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_13_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_13_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_13_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_13_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_13_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_13_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_13_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_13_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_13_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_13_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_13_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_14_clock; // @[Array.scala 41:54]
  wire  array_14_reset; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_14_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_14_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_14_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_14_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_14_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_14_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_14_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_14_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_14_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_14_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_14_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_14_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_14_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_14_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_14_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_14_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_14_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_14_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_14_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_14_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_14_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_14_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_14_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_14_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  wire  array_15_clock; // @[Array.scala 41:54]
  wire  array_15_reset; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_0_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_0_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_1_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_1_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_2_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_2_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_3_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_3_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_4_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_4_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_5_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_5_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_6_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_6_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_7_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_7_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_8_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_8_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_9_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_9_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_10_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_10_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_11_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_11_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_12_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_12_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_13_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_13_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_14_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_14_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_15_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_15_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_16_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_16_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_17_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_17_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_18_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_18_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_19_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_19_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_20_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_20_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_21_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_21_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_22_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_22_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_23_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_23_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_24_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_24_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_25_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_25_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_26_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_26_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_27_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_27_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_28_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_28_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_29_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_29_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_30_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_30_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_31_a; // @[Array.scala 41:54]
  wire  array_15_io_d_in_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_in_31_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_0_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_0_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_0_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_0_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_1_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_1_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_1_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_1_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_2_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_2_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_2_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_2_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_3_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_3_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_3_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_3_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_4_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_4_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_4_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_4_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_5_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_5_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_5_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_5_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_6_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_6_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_6_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_6_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_7_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_7_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_7_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_7_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_8_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_8_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_8_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_8_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_9_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_9_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_9_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_9_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_10_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_10_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_10_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_10_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_11_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_11_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_11_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_11_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_12_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_12_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_12_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_12_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_13_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_13_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_13_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_13_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_14_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_14_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_14_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_14_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_15_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_15_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_15_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_15_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_16_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_16_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_16_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_16_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_17_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_17_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_17_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_17_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_18_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_18_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_18_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_18_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_19_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_19_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_19_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_19_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_20_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_20_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_20_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_20_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_21_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_21_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_21_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_21_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_22_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_22_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_22_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_22_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_23_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_23_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_23_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_23_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_24_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_24_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_24_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_24_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_25_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_25_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_25_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_25_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_26_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_26_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_26_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_26_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_27_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_27_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_27_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_27_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_28_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_28_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_28_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_28_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_29_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_29_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_29_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_29_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_30_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_30_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_30_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_30_valid_b; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_31_a; // @[Array.scala 41:54]
  wire  array_15_io_d_out_31_valid_a; // @[Array.scala 41:54]
  wire [63:0] array_15_io_d_out_31_b; // @[Array.scala 41:54]
  wire  array_15_io_d_out_31_valid_b; // @[Array.scala 41:54]
  wire  array_15_io_wr_en_mem1; // @[Array.scala 41:54]
  wire  array_15_io_wr_en_mem2; // @[Array.scala 41:54]
  wire  array_15_io_wr_en_mem3; // @[Array.scala 41:54]
  wire  array_15_io_wr_en_mem4; // @[Array.scala 41:54]
  wire  array_15_io_wr_en_mem5; // @[Array.scala 41:54]
  wire  array_15_io_wr_en_mem6; // @[Array.scala 41:54]
  wire [287:0] array_15_io_wr_instr_mem1; // @[Array.scala 41:54]
  wire [127:0] array_15_io_wr_instr_mem2; // @[Array.scala 41:54]
  wire [127:0] array_15_io_wr_instr_mem3; // @[Array.scala 41:54]
  wire [127:0] array_15_io_wr_instr_mem4; // @[Array.scala 41:54]
  wire [127:0] array_15_io_wr_instr_mem5; // @[Array.scala 41:54]
  wire [127:0] array_15_io_wr_instr_mem6; // @[Array.scala 41:54]
  wire [7:0] array_15_io_PC1_in; // @[Array.scala 41:54]
  wire [7:0] array_15_io_PC6_out; // @[Array.scala 41:54]
  wire [7:0] array_15_io_Addr_in; // @[Array.scala 41:54]
  wire [7:0] array_15_io_Addr_out; // @[Array.scala 41:54]
  wire [1:0] array_15_io_Tag_in_Tag; // @[Array.scala 41:54]
  wire [2:0] array_15_io_Tag_in_RoundCnt; // @[Array.scala 41:54]
  wire [1:0] array_15_io_Tag_out_Tag; // @[Array.scala 41:54]
  wire [2:0] array_15_io_Tag_out_RoundCnt; // @[Array.scala 41:54]
  BuildingBlockNew array_0 ( // @[Array.scala 41:54]
    .clock(array_0_clock),
    .reset(array_0_reset),
    .io_d_in_0_a(array_0_io_d_in_0_a),
    .io_d_in_0_valid_a(array_0_io_d_in_0_valid_a),
    .io_d_in_0_b(array_0_io_d_in_0_b),
    .io_d_in_1_a(array_0_io_d_in_1_a),
    .io_d_in_1_valid_a(array_0_io_d_in_1_valid_a),
    .io_d_in_1_b(array_0_io_d_in_1_b),
    .io_d_in_2_a(array_0_io_d_in_2_a),
    .io_d_in_2_valid_a(array_0_io_d_in_2_valid_a),
    .io_d_in_2_b(array_0_io_d_in_2_b),
    .io_d_in_3_a(array_0_io_d_in_3_a),
    .io_d_in_3_valid_a(array_0_io_d_in_3_valid_a),
    .io_d_in_3_b(array_0_io_d_in_3_b),
    .io_d_in_4_a(array_0_io_d_in_4_a),
    .io_d_in_4_valid_a(array_0_io_d_in_4_valid_a),
    .io_d_in_4_b(array_0_io_d_in_4_b),
    .io_d_in_5_a(array_0_io_d_in_5_a),
    .io_d_in_5_valid_a(array_0_io_d_in_5_valid_a),
    .io_d_in_5_b(array_0_io_d_in_5_b),
    .io_d_in_6_a(array_0_io_d_in_6_a),
    .io_d_in_6_valid_a(array_0_io_d_in_6_valid_a),
    .io_d_in_6_b(array_0_io_d_in_6_b),
    .io_d_in_7_a(array_0_io_d_in_7_a),
    .io_d_in_7_valid_a(array_0_io_d_in_7_valid_a),
    .io_d_in_7_b(array_0_io_d_in_7_b),
    .io_d_in_8_a(array_0_io_d_in_8_a),
    .io_d_in_8_valid_a(array_0_io_d_in_8_valid_a),
    .io_d_in_8_b(array_0_io_d_in_8_b),
    .io_d_in_9_a(array_0_io_d_in_9_a),
    .io_d_in_9_valid_a(array_0_io_d_in_9_valid_a),
    .io_d_in_9_b(array_0_io_d_in_9_b),
    .io_d_in_10_a(array_0_io_d_in_10_a),
    .io_d_in_10_valid_a(array_0_io_d_in_10_valid_a),
    .io_d_in_10_b(array_0_io_d_in_10_b),
    .io_d_in_11_a(array_0_io_d_in_11_a),
    .io_d_in_11_valid_a(array_0_io_d_in_11_valid_a),
    .io_d_in_11_b(array_0_io_d_in_11_b),
    .io_d_in_12_a(array_0_io_d_in_12_a),
    .io_d_in_12_valid_a(array_0_io_d_in_12_valid_a),
    .io_d_in_12_b(array_0_io_d_in_12_b),
    .io_d_in_13_a(array_0_io_d_in_13_a),
    .io_d_in_13_valid_a(array_0_io_d_in_13_valid_a),
    .io_d_in_13_b(array_0_io_d_in_13_b),
    .io_d_in_14_a(array_0_io_d_in_14_a),
    .io_d_in_14_valid_a(array_0_io_d_in_14_valid_a),
    .io_d_in_14_b(array_0_io_d_in_14_b),
    .io_d_in_15_a(array_0_io_d_in_15_a),
    .io_d_in_15_valid_a(array_0_io_d_in_15_valid_a),
    .io_d_in_15_b(array_0_io_d_in_15_b),
    .io_d_in_16_a(array_0_io_d_in_16_a),
    .io_d_in_16_valid_a(array_0_io_d_in_16_valid_a),
    .io_d_in_16_b(array_0_io_d_in_16_b),
    .io_d_in_17_a(array_0_io_d_in_17_a),
    .io_d_in_17_valid_a(array_0_io_d_in_17_valid_a),
    .io_d_in_17_b(array_0_io_d_in_17_b),
    .io_d_in_18_a(array_0_io_d_in_18_a),
    .io_d_in_18_valid_a(array_0_io_d_in_18_valid_a),
    .io_d_in_18_b(array_0_io_d_in_18_b),
    .io_d_in_19_a(array_0_io_d_in_19_a),
    .io_d_in_19_valid_a(array_0_io_d_in_19_valid_a),
    .io_d_in_19_b(array_0_io_d_in_19_b),
    .io_d_in_20_a(array_0_io_d_in_20_a),
    .io_d_in_20_valid_a(array_0_io_d_in_20_valid_a),
    .io_d_in_20_b(array_0_io_d_in_20_b),
    .io_d_in_21_a(array_0_io_d_in_21_a),
    .io_d_in_21_valid_a(array_0_io_d_in_21_valid_a),
    .io_d_in_21_b(array_0_io_d_in_21_b),
    .io_d_in_22_a(array_0_io_d_in_22_a),
    .io_d_in_22_valid_a(array_0_io_d_in_22_valid_a),
    .io_d_in_22_b(array_0_io_d_in_22_b),
    .io_d_in_23_a(array_0_io_d_in_23_a),
    .io_d_in_23_valid_a(array_0_io_d_in_23_valid_a),
    .io_d_in_23_b(array_0_io_d_in_23_b),
    .io_d_in_24_a(array_0_io_d_in_24_a),
    .io_d_in_24_valid_a(array_0_io_d_in_24_valid_a),
    .io_d_in_24_b(array_0_io_d_in_24_b),
    .io_d_in_25_a(array_0_io_d_in_25_a),
    .io_d_in_25_valid_a(array_0_io_d_in_25_valid_a),
    .io_d_in_25_b(array_0_io_d_in_25_b),
    .io_d_in_26_a(array_0_io_d_in_26_a),
    .io_d_in_26_valid_a(array_0_io_d_in_26_valid_a),
    .io_d_in_26_b(array_0_io_d_in_26_b),
    .io_d_in_27_a(array_0_io_d_in_27_a),
    .io_d_in_27_valid_a(array_0_io_d_in_27_valid_a),
    .io_d_in_27_b(array_0_io_d_in_27_b),
    .io_d_in_28_a(array_0_io_d_in_28_a),
    .io_d_in_28_valid_a(array_0_io_d_in_28_valid_a),
    .io_d_in_28_b(array_0_io_d_in_28_b),
    .io_d_in_29_a(array_0_io_d_in_29_a),
    .io_d_in_29_valid_a(array_0_io_d_in_29_valid_a),
    .io_d_in_29_b(array_0_io_d_in_29_b),
    .io_d_in_30_a(array_0_io_d_in_30_a),
    .io_d_in_30_valid_a(array_0_io_d_in_30_valid_a),
    .io_d_in_30_b(array_0_io_d_in_30_b),
    .io_d_in_31_a(array_0_io_d_in_31_a),
    .io_d_in_31_valid_a(array_0_io_d_in_31_valid_a),
    .io_d_in_31_b(array_0_io_d_in_31_b),
    .io_d_out_0_a(array_0_io_d_out_0_a),
    .io_d_out_0_valid_a(array_0_io_d_out_0_valid_a),
    .io_d_out_0_b(array_0_io_d_out_0_b),
    .io_d_out_0_valid_b(array_0_io_d_out_0_valid_b),
    .io_d_out_1_a(array_0_io_d_out_1_a),
    .io_d_out_1_valid_a(array_0_io_d_out_1_valid_a),
    .io_d_out_1_b(array_0_io_d_out_1_b),
    .io_d_out_1_valid_b(array_0_io_d_out_1_valid_b),
    .io_d_out_2_a(array_0_io_d_out_2_a),
    .io_d_out_2_valid_a(array_0_io_d_out_2_valid_a),
    .io_d_out_2_b(array_0_io_d_out_2_b),
    .io_d_out_2_valid_b(array_0_io_d_out_2_valid_b),
    .io_d_out_3_a(array_0_io_d_out_3_a),
    .io_d_out_3_valid_a(array_0_io_d_out_3_valid_a),
    .io_d_out_3_b(array_0_io_d_out_3_b),
    .io_d_out_3_valid_b(array_0_io_d_out_3_valid_b),
    .io_d_out_4_a(array_0_io_d_out_4_a),
    .io_d_out_4_valid_a(array_0_io_d_out_4_valid_a),
    .io_d_out_4_b(array_0_io_d_out_4_b),
    .io_d_out_4_valid_b(array_0_io_d_out_4_valid_b),
    .io_d_out_5_a(array_0_io_d_out_5_a),
    .io_d_out_5_valid_a(array_0_io_d_out_5_valid_a),
    .io_d_out_5_b(array_0_io_d_out_5_b),
    .io_d_out_5_valid_b(array_0_io_d_out_5_valid_b),
    .io_d_out_6_a(array_0_io_d_out_6_a),
    .io_d_out_6_valid_a(array_0_io_d_out_6_valid_a),
    .io_d_out_6_b(array_0_io_d_out_6_b),
    .io_d_out_6_valid_b(array_0_io_d_out_6_valid_b),
    .io_d_out_7_a(array_0_io_d_out_7_a),
    .io_d_out_7_valid_a(array_0_io_d_out_7_valid_a),
    .io_d_out_7_b(array_0_io_d_out_7_b),
    .io_d_out_7_valid_b(array_0_io_d_out_7_valid_b),
    .io_d_out_8_a(array_0_io_d_out_8_a),
    .io_d_out_8_valid_a(array_0_io_d_out_8_valid_a),
    .io_d_out_8_b(array_0_io_d_out_8_b),
    .io_d_out_8_valid_b(array_0_io_d_out_8_valid_b),
    .io_d_out_9_a(array_0_io_d_out_9_a),
    .io_d_out_9_valid_a(array_0_io_d_out_9_valid_a),
    .io_d_out_9_b(array_0_io_d_out_9_b),
    .io_d_out_9_valid_b(array_0_io_d_out_9_valid_b),
    .io_d_out_10_a(array_0_io_d_out_10_a),
    .io_d_out_10_valid_a(array_0_io_d_out_10_valid_a),
    .io_d_out_10_b(array_0_io_d_out_10_b),
    .io_d_out_10_valid_b(array_0_io_d_out_10_valid_b),
    .io_d_out_11_a(array_0_io_d_out_11_a),
    .io_d_out_11_valid_a(array_0_io_d_out_11_valid_a),
    .io_d_out_11_b(array_0_io_d_out_11_b),
    .io_d_out_11_valid_b(array_0_io_d_out_11_valid_b),
    .io_d_out_12_a(array_0_io_d_out_12_a),
    .io_d_out_12_valid_a(array_0_io_d_out_12_valid_a),
    .io_d_out_12_b(array_0_io_d_out_12_b),
    .io_d_out_12_valid_b(array_0_io_d_out_12_valid_b),
    .io_d_out_13_a(array_0_io_d_out_13_a),
    .io_d_out_13_valid_a(array_0_io_d_out_13_valid_a),
    .io_d_out_13_b(array_0_io_d_out_13_b),
    .io_d_out_13_valid_b(array_0_io_d_out_13_valid_b),
    .io_d_out_14_a(array_0_io_d_out_14_a),
    .io_d_out_14_valid_a(array_0_io_d_out_14_valid_a),
    .io_d_out_14_b(array_0_io_d_out_14_b),
    .io_d_out_14_valid_b(array_0_io_d_out_14_valid_b),
    .io_d_out_15_a(array_0_io_d_out_15_a),
    .io_d_out_15_valid_a(array_0_io_d_out_15_valid_a),
    .io_d_out_15_b(array_0_io_d_out_15_b),
    .io_d_out_15_valid_b(array_0_io_d_out_15_valid_b),
    .io_d_out_16_a(array_0_io_d_out_16_a),
    .io_d_out_16_valid_a(array_0_io_d_out_16_valid_a),
    .io_d_out_16_b(array_0_io_d_out_16_b),
    .io_d_out_16_valid_b(array_0_io_d_out_16_valid_b),
    .io_d_out_17_a(array_0_io_d_out_17_a),
    .io_d_out_17_valid_a(array_0_io_d_out_17_valid_a),
    .io_d_out_17_b(array_0_io_d_out_17_b),
    .io_d_out_17_valid_b(array_0_io_d_out_17_valid_b),
    .io_d_out_18_a(array_0_io_d_out_18_a),
    .io_d_out_18_valid_a(array_0_io_d_out_18_valid_a),
    .io_d_out_18_b(array_0_io_d_out_18_b),
    .io_d_out_18_valid_b(array_0_io_d_out_18_valid_b),
    .io_d_out_19_a(array_0_io_d_out_19_a),
    .io_d_out_19_valid_a(array_0_io_d_out_19_valid_a),
    .io_d_out_19_b(array_0_io_d_out_19_b),
    .io_d_out_19_valid_b(array_0_io_d_out_19_valid_b),
    .io_d_out_20_a(array_0_io_d_out_20_a),
    .io_d_out_20_valid_a(array_0_io_d_out_20_valid_a),
    .io_d_out_20_b(array_0_io_d_out_20_b),
    .io_d_out_20_valid_b(array_0_io_d_out_20_valid_b),
    .io_d_out_21_a(array_0_io_d_out_21_a),
    .io_d_out_21_valid_a(array_0_io_d_out_21_valid_a),
    .io_d_out_21_b(array_0_io_d_out_21_b),
    .io_d_out_21_valid_b(array_0_io_d_out_21_valid_b),
    .io_d_out_22_a(array_0_io_d_out_22_a),
    .io_d_out_22_valid_a(array_0_io_d_out_22_valid_a),
    .io_d_out_22_b(array_0_io_d_out_22_b),
    .io_d_out_22_valid_b(array_0_io_d_out_22_valid_b),
    .io_d_out_23_a(array_0_io_d_out_23_a),
    .io_d_out_23_valid_a(array_0_io_d_out_23_valid_a),
    .io_d_out_23_b(array_0_io_d_out_23_b),
    .io_d_out_23_valid_b(array_0_io_d_out_23_valid_b),
    .io_d_out_24_a(array_0_io_d_out_24_a),
    .io_d_out_24_valid_a(array_0_io_d_out_24_valid_a),
    .io_d_out_24_b(array_0_io_d_out_24_b),
    .io_d_out_24_valid_b(array_0_io_d_out_24_valid_b),
    .io_d_out_25_a(array_0_io_d_out_25_a),
    .io_d_out_25_valid_a(array_0_io_d_out_25_valid_a),
    .io_d_out_25_b(array_0_io_d_out_25_b),
    .io_d_out_25_valid_b(array_0_io_d_out_25_valid_b),
    .io_d_out_26_a(array_0_io_d_out_26_a),
    .io_d_out_26_valid_a(array_0_io_d_out_26_valid_a),
    .io_d_out_26_b(array_0_io_d_out_26_b),
    .io_d_out_26_valid_b(array_0_io_d_out_26_valid_b),
    .io_d_out_27_a(array_0_io_d_out_27_a),
    .io_d_out_27_valid_a(array_0_io_d_out_27_valid_a),
    .io_d_out_27_b(array_0_io_d_out_27_b),
    .io_d_out_27_valid_b(array_0_io_d_out_27_valid_b),
    .io_d_out_28_a(array_0_io_d_out_28_a),
    .io_d_out_28_valid_a(array_0_io_d_out_28_valid_a),
    .io_d_out_28_b(array_0_io_d_out_28_b),
    .io_d_out_28_valid_b(array_0_io_d_out_28_valid_b),
    .io_d_out_29_a(array_0_io_d_out_29_a),
    .io_d_out_29_valid_a(array_0_io_d_out_29_valid_a),
    .io_d_out_29_b(array_0_io_d_out_29_b),
    .io_d_out_29_valid_b(array_0_io_d_out_29_valid_b),
    .io_d_out_30_a(array_0_io_d_out_30_a),
    .io_d_out_30_valid_a(array_0_io_d_out_30_valid_a),
    .io_d_out_30_b(array_0_io_d_out_30_b),
    .io_d_out_30_valid_b(array_0_io_d_out_30_valid_b),
    .io_d_out_31_a(array_0_io_d_out_31_a),
    .io_d_out_31_valid_a(array_0_io_d_out_31_valid_a),
    .io_d_out_31_b(array_0_io_d_out_31_b),
    .io_d_out_31_valid_b(array_0_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_0_io_wr_en_mem1),
    .io_wr_en_mem2(array_0_io_wr_en_mem2),
    .io_wr_en_mem3(array_0_io_wr_en_mem3),
    .io_wr_en_mem4(array_0_io_wr_en_mem4),
    .io_wr_en_mem5(array_0_io_wr_en_mem5),
    .io_wr_en_mem6(array_0_io_wr_en_mem6),
    .io_wr_instr_mem1(array_0_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_0_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_0_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_0_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_0_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_0_io_wr_instr_mem6),
    .io_PC1_in(array_0_io_PC1_in),
    .io_PC6_out(array_0_io_PC6_out),
    .io_Addr_in(array_0_io_Addr_in),
    .io_Addr_out(array_0_io_Addr_out),
    .io_Tag_in_Tag(array_0_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_0_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_0_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_0_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_1 ( // @[Array.scala 41:54]
    .clock(array_1_clock),
    .reset(array_1_reset),
    .io_d_in_0_a(array_1_io_d_in_0_a),
    .io_d_in_0_valid_a(array_1_io_d_in_0_valid_a),
    .io_d_in_0_b(array_1_io_d_in_0_b),
    .io_d_in_1_a(array_1_io_d_in_1_a),
    .io_d_in_1_valid_a(array_1_io_d_in_1_valid_a),
    .io_d_in_1_b(array_1_io_d_in_1_b),
    .io_d_in_2_a(array_1_io_d_in_2_a),
    .io_d_in_2_valid_a(array_1_io_d_in_2_valid_a),
    .io_d_in_2_b(array_1_io_d_in_2_b),
    .io_d_in_3_a(array_1_io_d_in_3_a),
    .io_d_in_3_valid_a(array_1_io_d_in_3_valid_a),
    .io_d_in_3_b(array_1_io_d_in_3_b),
    .io_d_in_4_a(array_1_io_d_in_4_a),
    .io_d_in_4_valid_a(array_1_io_d_in_4_valid_a),
    .io_d_in_4_b(array_1_io_d_in_4_b),
    .io_d_in_5_a(array_1_io_d_in_5_a),
    .io_d_in_5_valid_a(array_1_io_d_in_5_valid_a),
    .io_d_in_5_b(array_1_io_d_in_5_b),
    .io_d_in_6_a(array_1_io_d_in_6_a),
    .io_d_in_6_valid_a(array_1_io_d_in_6_valid_a),
    .io_d_in_6_b(array_1_io_d_in_6_b),
    .io_d_in_7_a(array_1_io_d_in_7_a),
    .io_d_in_7_valid_a(array_1_io_d_in_7_valid_a),
    .io_d_in_7_b(array_1_io_d_in_7_b),
    .io_d_in_8_a(array_1_io_d_in_8_a),
    .io_d_in_8_valid_a(array_1_io_d_in_8_valid_a),
    .io_d_in_8_b(array_1_io_d_in_8_b),
    .io_d_in_9_a(array_1_io_d_in_9_a),
    .io_d_in_9_valid_a(array_1_io_d_in_9_valid_a),
    .io_d_in_9_b(array_1_io_d_in_9_b),
    .io_d_in_10_a(array_1_io_d_in_10_a),
    .io_d_in_10_valid_a(array_1_io_d_in_10_valid_a),
    .io_d_in_10_b(array_1_io_d_in_10_b),
    .io_d_in_11_a(array_1_io_d_in_11_a),
    .io_d_in_11_valid_a(array_1_io_d_in_11_valid_a),
    .io_d_in_11_b(array_1_io_d_in_11_b),
    .io_d_in_12_a(array_1_io_d_in_12_a),
    .io_d_in_12_valid_a(array_1_io_d_in_12_valid_a),
    .io_d_in_12_b(array_1_io_d_in_12_b),
    .io_d_in_13_a(array_1_io_d_in_13_a),
    .io_d_in_13_valid_a(array_1_io_d_in_13_valid_a),
    .io_d_in_13_b(array_1_io_d_in_13_b),
    .io_d_in_14_a(array_1_io_d_in_14_a),
    .io_d_in_14_valid_a(array_1_io_d_in_14_valid_a),
    .io_d_in_14_b(array_1_io_d_in_14_b),
    .io_d_in_15_a(array_1_io_d_in_15_a),
    .io_d_in_15_valid_a(array_1_io_d_in_15_valid_a),
    .io_d_in_15_b(array_1_io_d_in_15_b),
    .io_d_in_16_a(array_1_io_d_in_16_a),
    .io_d_in_16_valid_a(array_1_io_d_in_16_valid_a),
    .io_d_in_16_b(array_1_io_d_in_16_b),
    .io_d_in_17_a(array_1_io_d_in_17_a),
    .io_d_in_17_valid_a(array_1_io_d_in_17_valid_a),
    .io_d_in_17_b(array_1_io_d_in_17_b),
    .io_d_in_18_a(array_1_io_d_in_18_a),
    .io_d_in_18_valid_a(array_1_io_d_in_18_valid_a),
    .io_d_in_18_b(array_1_io_d_in_18_b),
    .io_d_in_19_a(array_1_io_d_in_19_a),
    .io_d_in_19_valid_a(array_1_io_d_in_19_valid_a),
    .io_d_in_19_b(array_1_io_d_in_19_b),
    .io_d_in_20_a(array_1_io_d_in_20_a),
    .io_d_in_20_valid_a(array_1_io_d_in_20_valid_a),
    .io_d_in_20_b(array_1_io_d_in_20_b),
    .io_d_in_21_a(array_1_io_d_in_21_a),
    .io_d_in_21_valid_a(array_1_io_d_in_21_valid_a),
    .io_d_in_21_b(array_1_io_d_in_21_b),
    .io_d_in_22_a(array_1_io_d_in_22_a),
    .io_d_in_22_valid_a(array_1_io_d_in_22_valid_a),
    .io_d_in_22_b(array_1_io_d_in_22_b),
    .io_d_in_23_a(array_1_io_d_in_23_a),
    .io_d_in_23_valid_a(array_1_io_d_in_23_valid_a),
    .io_d_in_23_b(array_1_io_d_in_23_b),
    .io_d_in_24_a(array_1_io_d_in_24_a),
    .io_d_in_24_valid_a(array_1_io_d_in_24_valid_a),
    .io_d_in_24_b(array_1_io_d_in_24_b),
    .io_d_in_25_a(array_1_io_d_in_25_a),
    .io_d_in_25_valid_a(array_1_io_d_in_25_valid_a),
    .io_d_in_25_b(array_1_io_d_in_25_b),
    .io_d_in_26_a(array_1_io_d_in_26_a),
    .io_d_in_26_valid_a(array_1_io_d_in_26_valid_a),
    .io_d_in_26_b(array_1_io_d_in_26_b),
    .io_d_in_27_a(array_1_io_d_in_27_a),
    .io_d_in_27_valid_a(array_1_io_d_in_27_valid_a),
    .io_d_in_27_b(array_1_io_d_in_27_b),
    .io_d_in_28_a(array_1_io_d_in_28_a),
    .io_d_in_28_valid_a(array_1_io_d_in_28_valid_a),
    .io_d_in_28_b(array_1_io_d_in_28_b),
    .io_d_in_29_a(array_1_io_d_in_29_a),
    .io_d_in_29_valid_a(array_1_io_d_in_29_valid_a),
    .io_d_in_29_b(array_1_io_d_in_29_b),
    .io_d_in_30_a(array_1_io_d_in_30_a),
    .io_d_in_30_valid_a(array_1_io_d_in_30_valid_a),
    .io_d_in_30_b(array_1_io_d_in_30_b),
    .io_d_in_31_a(array_1_io_d_in_31_a),
    .io_d_in_31_valid_a(array_1_io_d_in_31_valid_a),
    .io_d_in_31_b(array_1_io_d_in_31_b),
    .io_d_out_0_a(array_1_io_d_out_0_a),
    .io_d_out_0_valid_a(array_1_io_d_out_0_valid_a),
    .io_d_out_0_b(array_1_io_d_out_0_b),
    .io_d_out_0_valid_b(array_1_io_d_out_0_valid_b),
    .io_d_out_1_a(array_1_io_d_out_1_a),
    .io_d_out_1_valid_a(array_1_io_d_out_1_valid_a),
    .io_d_out_1_b(array_1_io_d_out_1_b),
    .io_d_out_1_valid_b(array_1_io_d_out_1_valid_b),
    .io_d_out_2_a(array_1_io_d_out_2_a),
    .io_d_out_2_valid_a(array_1_io_d_out_2_valid_a),
    .io_d_out_2_b(array_1_io_d_out_2_b),
    .io_d_out_2_valid_b(array_1_io_d_out_2_valid_b),
    .io_d_out_3_a(array_1_io_d_out_3_a),
    .io_d_out_3_valid_a(array_1_io_d_out_3_valid_a),
    .io_d_out_3_b(array_1_io_d_out_3_b),
    .io_d_out_3_valid_b(array_1_io_d_out_3_valid_b),
    .io_d_out_4_a(array_1_io_d_out_4_a),
    .io_d_out_4_valid_a(array_1_io_d_out_4_valid_a),
    .io_d_out_4_b(array_1_io_d_out_4_b),
    .io_d_out_4_valid_b(array_1_io_d_out_4_valid_b),
    .io_d_out_5_a(array_1_io_d_out_5_a),
    .io_d_out_5_valid_a(array_1_io_d_out_5_valid_a),
    .io_d_out_5_b(array_1_io_d_out_5_b),
    .io_d_out_5_valid_b(array_1_io_d_out_5_valid_b),
    .io_d_out_6_a(array_1_io_d_out_6_a),
    .io_d_out_6_valid_a(array_1_io_d_out_6_valid_a),
    .io_d_out_6_b(array_1_io_d_out_6_b),
    .io_d_out_6_valid_b(array_1_io_d_out_6_valid_b),
    .io_d_out_7_a(array_1_io_d_out_7_a),
    .io_d_out_7_valid_a(array_1_io_d_out_7_valid_a),
    .io_d_out_7_b(array_1_io_d_out_7_b),
    .io_d_out_7_valid_b(array_1_io_d_out_7_valid_b),
    .io_d_out_8_a(array_1_io_d_out_8_a),
    .io_d_out_8_valid_a(array_1_io_d_out_8_valid_a),
    .io_d_out_8_b(array_1_io_d_out_8_b),
    .io_d_out_8_valid_b(array_1_io_d_out_8_valid_b),
    .io_d_out_9_a(array_1_io_d_out_9_a),
    .io_d_out_9_valid_a(array_1_io_d_out_9_valid_a),
    .io_d_out_9_b(array_1_io_d_out_9_b),
    .io_d_out_9_valid_b(array_1_io_d_out_9_valid_b),
    .io_d_out_10_a(array_1_io_d_out_10_a),
    .io_d_out_10_valid_a(array_1_io_d_out_10_valid_a),
    .io_d_out_10_b(array_1_io_d_out_10_b),
    .io_d_out_10_valid_b(array_1_io_d_out_10_valid_b),
    .io_d_out_11_a(array_1_io_d_out_11_a),
    .io_d_out_11_valid_a(array_1_io_d_out_11_valid_a),
    .io_d_out_11_b(array_1_io_d_out_11_b),
    .io_d_out_11_valid_b(array_1_io_d_out_11_valid_b),
    .io_d_out_12_a(array_1_io_d_out_12_a),
    .io_d_out_12_valid_a(array_1_io_d_out_12_valid_a),
    .io_d_out_12_b(array_1_io_d_out_12_b),
    .io_d_out_12_valid_b(array_1_io_d_out_12_valid_b),
    .io_d_out_13_a(array_1_io_d_out_13_a),
    .io_d_out_13_valid_a(array_1_io_d_out_13_valid_a),
    .io_d_out_13_b(array_1_io_d_out_13_b),
    .io_d_out_13_valid_b(array_1_io_d_out_13_valid_b),
    .io_d_out_14_a(array_1_io_d_out_14_a),
    .io_d_out_14_valid_a(array_1_io_d_out_14_valid_a),
    .io_d_out_14_b(array_1_io_d_out_14_b),
    .io_d_out_14_valid_b(array_1_io_d_out_14_valid_b),
    .io_d_out_15_a(array_1_io_d_out_15_a),
    .io_d_out_15_valid_a(array_1_io_d_out_15_valid_a),
    .io_d_out_15_b(array_1_io_d_out_15_b),
    .io_d_out_15_valid_b(array_1_io_d_out_15_valid_b),
    .io_d_out_16_a(array_1_io_d_out_16_a),
    .io_d_out_16_valid_a(array_1_io_d_out_16_valid_a),
    .io_d_out_16_b(array_1_io_d_out_16_b),
    .io_d_out_16_valid_b(array_1_io_d_out_16_valid_b),
    .io_d_out_17_a(array_1_io_d_out_17_a),
    .io_d_out_17_valid_a(array_1_io_d_out_17_valid_a),
    .io_d_out_17_b(array_1_io_d_out_17_b),
    .io_d_out_17_valid_b(array_1_io_d_out_17_valid_b),
    .io_d_out_18_a(array_1_io_d_out_18_a),
    .io_d_out_18_valid_a(array_1_io_d_out_18_valid_a),
    .io_d_out_18_b(array_1_io_d_out_18_b),
    .io_d_out_18_valid_b(array_1_io_d_out_18_valid_b),
    .io_d_out_19_a(array_1_io_d_out_19_a),
    .io_d_out_19_valid_a(array_1_io_d_out_19_valid_a),
    .io_d_out_19_b(array_1_io_d_out_19_b),
    .io_d_out_19_valid_b(array_1_io_d_out_19_valid_b),
    .io_d_out_20_a(array_1_io_d_out_20_a),
    .io_d_out_20_valid_a(array_1_io_d_out_20_valid_a),
    .io_d_out_20_b(array_1_io_d_out_20_b),
    .io_d_out_20_valid_b(array_1_io_d_out_20_valid_b),
    .io_d_out_21_a(array_1_io_d_out_21_a),
    .io_d_out_21_valid_a(array_1_io_d_out_21_valid_a),
    .io_d_out_21_b(array_1_io_d_out_21_b),
    .io_d_out_21_valid_b(array_1_io_d_out_21_valid_b),
    .io_d_out_22_a(array_1_io_d_out_22_a),
    .io_d_out_22_valid_a(array_1_io_d_out_22_valid_a),
    .io_d_out_22_b(array_1_io_d_out_22_b),
    .io_d_out_22_valid_b(array_1_io_d_out_22_valid_b),
    .io_d_out_23_a(array_1_io_d_out_23_a),
    .io_d_out_23_valid_a(array_1_io_d_out_23_valid_a),
    .io_d_out_23_b(array_1_io_d_out_23_b),
    .io_d_out_23_valid_b(array_1_io_d_out_23_valid_b),
    .io_d_out_24_a(array_1_io_d_out_24_a),
    .io_d_out_24_valid_a(array_1_io_d_out_24_valid_a),
    .io_d_out_24_b(array_1_io_d_out_24_b),
    .io_d_out_24_valid_b(array_1_io_d_out_24_valid_b),
    .io_d_out_25_a(array_1_io_d_out_25_a),
    .io_d_out_25_valid_a(array_1_io_d_out_25_valid_a),
    .io_d_out_25_b(array_1_io_d_out_25_b),
    .io_d_out_25_valid_b(array_1_io_d_out_25_valid_b),
    .io_d_out_26_a(array_1_io_d_out_26_a),
    .io_d_out_26_valid_a(array_1_io_d_out_26_valid_a),
    .io_d_out_26_b(array_1_io_d_out_26_b),
    .io_d_out_26_valid_b(array_1_io_d_out_26_valid_b),
    .io_d_out_27_a(array_1_io_d_out_27_a),
    .io_d_out_27_valid_a(array_1_io_d_out_27_valid_a),
    .io_d_out_27_b(array_1_io_d_out_27_b),
    .io_d_out_27_valid_b(array_1_io_d_out_27_valid_b),
    .io_d_out_28_a(array_1_io_d_out_28_a),
    .io_d_out_28_valid_a(array_1_io_d_out_28_valid_a),
    .io_d_out_28_b(array_1_io_d_out_28_b),
    .io_d_out_28_valid_b(array_1_io_d_out_28_valid_b),
    .io_d_out_29_a(array_1_io_d_out_29_a),
    .io_d_out_29_valid_a(array_1_io_d_out_29_valid_a),
    .io_d_out_29_b(array_1_io_d_out_29_b),
    .io_d_out_29_valid_b(array_1_io_d_out_29_valid_b),
    .io_d_out_30_a(array_1_io_d_out_30_a),
    .io_d_out_30_valid_a(array_1_io_d_out_30_valid_a),
    .io_d_out_30_b(array_1_io_d_out_30_b),
    .io_d_out_30_valid_b(array_1_io_d_out_30_valid_b),
    .io_d_out_31_a(array_1_io_d_out_31_a),
    .io_d_out_31_valid_a(array_1_io_d_out_31_valid_a),
    .io_d_out_31_b(array_1_io_d_out_31_b),
    .io_d_out_31_valid_b(array_1_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_1_io_wr_en_mem1),
    .io_wr_en_mem2(array_1_io_wr_en_mem2),
    .io_wr_en_mem3(array_1_io_wr_en_mem3),
    .io_wr_en_mem4(array_1_io_wr_en_mem4),
    .io_wr_en_mem5(array_1_io_wr_en_mem5),
    .io_wr_en_mem6(array_1_io_wr_en_mem6),
    .io_wr_instr_mem1(array_1_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_1_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_1_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_1_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_1_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_1_io_wr_instr_mem6),
    .io_PC1_in(array_1_io_PC1_in),
    .io_PC6_out(array_1_io_PC6_out),
    .io_Addr_in(array_1_io_Addr_in),
    .io_Addr_out(array_1_io_Addr_out),
    .io_Tag_in_Tag(array_1_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_1_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_1_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_1_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_2 ( // @[Array.scala 41:54]
    .clock(array_2_clock),
    .reset(array_2_reset),
    .io_d_in_0_a(array_2_io_d_in_0_a),
    .io_d_in_0_valid_a(array_2_io_d_in_0_valid_a),
    .io_d_in_0_b(array_2_io_d_in_0_b),
    .io_d_in_1_a(array_2_io_d_in_1_a),
    .io_d_in_1_valid_a(array_2_io_d_in_1_valid_a),
    .io_d_in_1_b(array_2_io_d_in_1_b),
    .io_d_in_2_a(array_2_io_d_in_2_a),
    .io_d_in_2_valid_a(array_2_io_d_in_2_valid_a),
    .io_d_in_2_b(array_2_io_d_in_2_b),
    .io_d_in_3_a(array_2_io_d_in_3_a),
    .io_d_in_3_valid_a(array_2_io_d_in_3_valid_a),
    .io_d_in_3_b(array_2_io_d_in_3_b),
    .io_d_in_4_a(array_2_io_d_in_4_a),
    .io_d_in_4_valid_a(array_2_io_d_in_4_valid_a),
    .io_d_in_4_b(array_2_io_d_in_4_b),
    .io_d_in_5_a(array_2_io_d_in_5_a),
    .io_d_in_5_valid_a(array_2_io_d_in_5_valid_a),
    .io_d_in_5_b(array_2_io_d_in_5_b),
    .io_d_in_6_a(array_2_io_d_in_6_a),
    .io_d_in_6_valid_a(array_2_io_d_in_6_valid_a),
    .io_d_in_6_b(array_2_io_d_in_6_b),
    .io_d_in_7_a(array_2_io_d_in_7_a),
    .io_d_in_7_valid_a(array_2_io_d_in_7_valid_a),
    .io_d_in_7_b(array_2_io_d_in_7_b),
    .io_d_in_8_a(array_2_io_d_in_8_a),
    .io_d_in_8_valid_a(array_2_io_d_in_8_valid_a),
    .io_d_in_8_b(array_2_io_d_in_8_b),
    .io_d_in_9_a(array_2_io_d_in_9_a),
    .io_d_in_9_valid_a(array_2_io_d_in_9_valid_a),
    .io_d_in_9_b(array_2_io_d_in_9_b),
    .io_d_in_10_a(array_2_io_d_in_10_a),
    .io_d_in_10_valid_a(array_2_io_d_in_10_valid_a),
    .io_d_in_10_b(array_2_io_d_in_10_b),
    .io_d_in_11_a(array_2_io_d_in_11_a),
    .io_d_in_11_valid_a(array_2_io_d_in_11_valid_a),
    .io_d_in_11_b(array_2_io_d_in_11_b),
    .io_d_in_12_a(array_2_io_d_in_12_a),
    .io_d_in_12_valid_a(array_2_io_d_in_12_valid_a),
    .io_d_in_12_b(array_2_io_d_in_12_b),
    .io_d_in_13_a(array_2_io_d_in_13_a),
    .io_d_in_13_valid_a(array_2_io_d_in_13_valid_a),
    .io_d_in_13_b(array_2_io_d_in_13_b),
    .io_d_in_14_a(array_2_io_d_in_14_a),
    .io_d_in_14_valid_a(array_2_io_d_in_14_valid_a),
    .io_d_in_14_b(array_2_io_d_in_14_b),
    .io_d_in_15_a(array_2_io_d_in_15_a),
    .io_d_in_15_valid_a(array_2_io_d_in_15_valid_a),
    .io_d_in_15_b(array_2_io_d_in_15_b),
    .io_d_in_16_a(array_2_io_d_in_16_a),
    .io_d_in_16_valid_a(array_2_io_d_in_16_valid_a),
    .io_d_in_16_b(array_2_io_d_in_16_b),
    .io_d_in_17_a(array_2_io_d_in_17_a),
    .io_d_in_17_valid_a(array_2_io_d_in_17_valid_a),
    .io_d_in_17_b(array_2_io_d_in_17_b),
    .io_d_in_18_a(array_2_io_d_in_18_a),
    .io_d_in_18_valid_a(array_2_io_d_in_18_valid_a),
    .io_d_in_18_b(array_2_io_d_in_18_b),
    .io_d_in_19_a(array_2_io_d_in_19_a),
    .io_d_in_19_valid_a(array_2_io_d_in_19_valid_a),
    .io_d_in_19_b(array_2_io_d_in_19_b),
    .io_d_in_20_a(array_2_io_d_in_20_a),
    .io_d_in_20_valid_a(array_2_io_d_in_20_valid_a),
    .io_d_in_20_b(array_2_io_d_in_20_b),
    .io_d_in_21_a(array_2_io_d_in_21_a),
    .io_d_in_21_valid_a(array_2_io_d_in_21_valid_a),
    .io_d_in_21_b(array_2_io_d_in_21_b),
    .io_d_in_22_a(array_2_io_d_in_22_a),
    .io_d_in_22_valid_a(array_2_io_d_in_22_valid_a),
    .io_d_in_22_b(array_2_io_d_in_22_b),
    .io_d_in_23_a(array_2_io_d_in_23_a),
    .io_d_in_23_valid_a(array_2_io_d_in_23_valid_a),
    .io_d_in_23_b(array_2_io_d_in_23_b),
    .io_d_in_24_a(array_2_io_d_in_24_a),
    .io_d_in_24_valid_a(array_2_io_d_in_24_valid_a),
    .io_d_in_24_b(array_2_io_d_in_24_b),
    .io_d_in_25_a(array_2_io_d_in_25_a),
    .io_d_in_25_valid_a(array_2_io_d_in_25_valid_a),
    .io_d_in_25_b(array_2_io_d_in_25_b),
    .io_d_in_26_a(array_2_io_d_in_26_a),
    .io_d_in_26_valid_a(array_2_io_d_in_26_valid_a),
    .io_d_in_26_b(array_2_io_d_in_26_b),
    .io_d_in_27_a(array_2_io_d_in_27_a),
    .io_d_in_27_valid_a(array_2_io_d_in_27_valid_a),
    .io_d_in_27_b(array_2_io_d_in_27_b),
    .io_d_in_28_a(array_2_io_d_in_28_a),
    .io_d_in_28_valid_a(array_2_io_d_in_28_valid_a),
    .io_d_in_28_b(array_2_io_d_in_28_b),
    .io_d_in_29_a(array_2_io_d_in_29_a),
    .io_d_in_29_valid_a(array_2_io_d_in_29_valid_a),
    .io_d_in_29_b(array_2_io_d_in_29_b),
    .io_d_in_30_a(array_2_io_d_in_30_a),
    .io_d_in_30_valid_a(array_2_io_d_in_30_valid_a),
    .io_d_in_30_b(array_2_io_d_in_30_b),
    .io_d_in_31_a(array_2_io_d_in_31_a),
    .io_d_in_31_valid_a(array_2_io_d_in_31_valid_a),
    .io_d_in_31_b(array_2_io_d_in_31_b),
    .io_d_out_0_a(array_2_io_d_out_0_a),
    .io_d_out_0_valid_a(array_2_io_d_out_0_valid_a),
    .io_d_out_0_b(array_2_io_d_out_0_b),
    .io_d_out_0_valid_b(array_2_io_d_out_0_valid_b),
    .io_d_out_1_a(array_2_io_d_out_1_a),
    .io_d_out_1_valid_a(array_2_io_d_out_1_valid_a),
    .io_d_out_1_b(array_2_io_d_out_1_b),
    .io_d_out_1_valid_b(array_2_io_d_out_1_valid_b),
    .io_d_out_2_a(array_2_io_d_out_2_a),
    .io_d_out_2_valid_a(array_2_io_d_out_2_valid_a),
    .io_d_out_2_b(array_2_io_d_out_2_b),
    .io_d_out_2_valid_b(array_2_io_d_out_2_valid_b),
    .io_d_out_3_a(array_2_io_d_out_3_a),
    .io_d_out_3_valid_a(array_2_io_d_out_3_valid_a),
    .io_d_out_3_b(array_2_io_d_out_3_b),
    .io_d_out_3_valid_b(array_2_io_d_out_3_valid_b),
    .io_d_out_4_a(array_2_io_d_out_4_a),
    .io_d_out_4_valid_a(array_2_io_d_out_4_valid_a),
    .io_d_out_4_b(array_2_io_d_out_4_b),
    .io_d_out_4_valid_b(array_2_io_d_out_4_valid_b),
    .io_d_out_5_a(array_2_io_d_out_5_a),
    .io_d_out_5_valid_a(array_2_io_d_out_5_valid_a),
    .io_d_out_5_b(array_2_io_d_out_5_b),
    .io_d_out_5_valid_b(array_2_io_d_out_5_valid_b),
    .io_d_out_6_a(array_2_io_d_out_6_a),
    .io_d_out_6_valid_a(array_2_io_d_out_6_valid_a),
    .io_d_out_6_b(array_2_io_d_out_6_b),
    .io_d_out_6_valid_b(array_2_io_d_out_6_valid_b),
    .io_d_out_7_a(array_2_io_d_out_7_a),
    .io_d_out_7_valid_a(array_2_io_d_out_7_valid_a),
    .io_d_out_7_b(array_2_io_d_out_7_b),
    .io_d_out_7_valid_b(array_2_io_d_out_7_valid_b),
    .io_d_out_8_a(array_2_io_d_out_8_a),
    .io_d_out_8_valid_a(array_2_io_d_out_8_valid_a),
    .io_d_out_8_b(array_2_io_d_out_8_b),
    .io_d_out_8_valid_b(array_2_io_d_out_8_valid_b),
    .io_d_out_9_a(array_2_io_d_out_9_a),
    .io_d_out_9_valid_a(array_2_io_d_out_9_valid_a),
    .io_d_out_9_b(array_2_io_d_out_9_b),
    .io_d_out_9_valid_b(array_2_io_d_out_9_valid_b),
    .io_d_out_10_a(array_2_io_d_out_10_a),
    .io_d_out_10_valid_a(array_2_io_d_out_10_valid_a),
    .io_d_out_10_b(array_2_io_d_out_10_b),
    .io_d_out_10_valid_b(array_2_io_d_out_10_valid_b),
    .io_d_out_11_a(array_2_io_d_out_11_a),
    .io_d_out_11_valid_a(array_2_io_d_out_11_valid_a),
    .io_d_out_11_b(array_2_io_d_out_11_b),
    .io_d_out_11_valid_b(array_2_io_d_out_11_valid_b),
    .io_d_out_12_a(array_2_io_d_out_12_a),
    .io_d_out_12_valid_a(array_2_io_d_out_12_valid_a),
    .io_d_out_12_b(array_2_io_d_out_12_b),
    .io_d_out_12_valid_b(array_2_io_d_out_12_valid_b),
    .io_d_out_13_a(array_2_io_d_out_13_a),
    .io_d_out_13_valid_a(array_2_io_d_out_13_valid_a),
    .io_d_out_13_b(array_2_io_d_out_13_b),
    .io_d_out_13_valid_b(array_2_io_d_out_13_valid_b),
    .io_d_out_14_a(array_2_io_d_out_14_a),
    .io_d_out_14_valid_a(array_2_io_d_out_14_valid_a),
    .io_d_out_14_b(array_2_io_d_out_14_b),
    .io_d_out_14_valid_b(array_2_io_d_out_14_valid_b),
    .io_d_out_15_a(array_2_io_d_out_15_a),
    .io_d_out_15_valid_a(array_2_io_d_out_15_valid_a),
    .io_d_out_15_b(array_2_io_d_out_15_b),
    .io_d_out_15_valid_b(array_2_io_d_out_15_valid_b),
    .io_d_out_16_a(array_2_io_d_out_16_a),
    .io_d_out_16_valid_a(array_2_io_d_out_16_valid_a),
    .io_d_out_16_b(array_2_io_d_out_16_b),
    .io_d_out_16_valid_b(array_2_io_d_out_16_valid_b),
    .io_d_out_17_a(array_2_io_d_out_17_a),
    .io_d_out_17_valid_a(array_2_io_d_out_17_valid_a),
    .io_d_out_17_b(array_2_io_d_out_17_b),
    .io_d_out_17_valid_b(array_2_io_d_out_17_valid_b),
    .io_d_out_18_a(array_2_io_d_out_18_a),
    .io_d_out_18_valid_a(array_2_io_d_out_18_valid_a),
    .io_d_out_18_b(array_2_io_d_out_18_b),
    .io_d_out_18_valid_b(array_2_io_d_out_18_valid_b),
    .io_d_out_19_a(array_2_io_d_out_19_a),
    .io_d_out_19_valid_a(array_2_io_d_out_19_valid_a),
    .io_d_out_19_b(array_2_io_d_out_19_b),
    .io_d_out_19_valid_b(array_2_io_d_out_19_valid_b),
    .io_d_out_20_a(array_2_io_d_out_20_a),
    .io_d_out_20_valid_a(array_2_io_d_out_20_valid_a),
    .io_d_out_20_b(array_2_io_d_out_20_b),
    .io_d_out_20_valid_b(array_2_io_d_out_20_valid_b),
    .io_d_out_21_a(array_2_io_d_out_21_a),
    .io_d_out_21_valid_a(array_2_io_d_out_21_valid_a),
    .io_d_out_21_b(array_2_io_d_out_21_b),
    .io_d_out_21_valid_b(array_2_io_d_out_21_valid_b),
    .io_d_out_22_a(array_2_io_d_out_22_a),
    .io_d_out_22_valid_a(array_2_io_d_out_22_valid_a),
    .io_d_out_22_b(array_2_io_d_out_22_b),
    .io_d_out_22_valid_b(array_2_io_d_out_22_valid_b),
    .io_d_out_23_a(array_2_io_d_out_23_a),
    .io_d_out_23_valid_a(array_2_io_d_out_23_valid_a),
    .io_d_out_23_b(array_2_io_d_out_23_b),
    .io_d_out_23_valid_b(array_2_io_d_out_23_valid_b),
    .io_d_out_24_a(array_2_io_d_out_24_a),
    .io_d_out_24_valid_a(array_2_io_d_out_24_valid_a),
    .io_d_out_24_b(array_2_io_d_out_24_b),
    .io_d_out_24_valid_b(array_2_io_d_out_24_valid_b),
    .io_d_out_25_a(array_2_io_d_out_25_a),
    .io_d_out_25_valid_a(array_2_io_d_out_25_valid_a),
    .io_d_out_25_b(array_2_io_d_out_25_b),
    .io_d_out_25_valid_b(array_2_io_d_out_25_valid_b),
    .io_d_out_26_a(array_2_io_d_out_26_a),
    .io_d_out_26_valid_a(array_2_io_d_out_26_valid_a),
    .io_d_out_26_b(array_2_io_d_out_26_b),
    .io_d_out_26_valid_b(array_2_io_d_out_26_valid_b),
    .io_d_out_27_a(array_2_io_d_out_27_a),
    .io_d_out_27_valid_a(array_2_io_d_out_27_valid_a),
    .io_d_out_27_b(array_2_io_d_out_27_b),
    .io_d_out_27_valid_b(array_2_io_d_out_27_valid_b),
    .io_d_out_28_a(array_2_io_d_out_28_a),
    .io_d_out_28_valid_a(array_2_io_d_out_28_valid_a),
    .io_d_out_28_b(array_2_io_d_out_28_b),
    .io_d_out_28_valid_b(array_2_io_d_out_28_valid_b),
    .io_d_out_29_a(array_2_io_d_out_29_a),
    .io_d_out_29_valid_a(array_2_io_d_out_29_valid_a),
    .io_d_out_29_b(array_2_io_d_out_29_b),
    .io_d_out_29_valid_b(array_2_io_d_out_29_valid_b),
    .io_d_out_30_a(array_2_io_d_out_30_a),
    .io_d_out_30_valid_a(array_2_io_d_out_30_valid_a),
    .io_d_out_30_b(array_2_io_d_out_30_b),
    .io_d_out_30_valid_b(array_2_io_d_out_30_valid_b),
    .io_d_out_31_a(array_2_io_d_out_31_a),
    .io_d_out_31_valid_a(array_2_io_d_out_31_valid_a),
    .io_d_out_31_b(array_2_io_d_out_31_b),
    .io_d_out_31_valid_b(array_2_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_2_io_wr_en_mem1),
    .io_wr_en_mem2(array_2_io_wr_en_mem2),
    .io_wr_en_mem3(array_2_io_wr_en_mem3),
    .io_wr_en_mem4(array_2_io_wr_en_mem4),
    .io_wr_en_mem5(array_2_io_wr_en_mem5),
    .io_wr_en_mem6(array_2_io_wr_en_mem6),
    .io_wr_instr_mem1(array_2_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_2_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_2_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_2_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_2_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_2_io_wr_instr_mem6),
    .io_PC1_in(array_2_io_PC1_in),
    .io_PC6_out(array_2_io_PC6_out),
    .io_Addr_in(array_2_io_Addr_in),
    .io_Addr_out(array_2_io_Addr_out),
    .io_Tag_in_Tag(array_2_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_2_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_2_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_2_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_3 ( // @[Array.scala 41:54]
    .clock(array_3_clock),
    .reset(array_3_reset),
    .io_d_in_0_a(array_3_io_d_in_0_a),
    .io_d_in_0_valid_a(array_3_io_d_in_0_valid_a),
    .io_d_in_0_b(array_3_io_d_in_0_b),
    .io_d_in_1_a(array_3_io_d_in_1_a),
    .io_d_in_1_valid_a(array_3_io_d_in_1_valid_a),
    .io_d_in_1_b(array_3_io_d_in_1_b),
    .io_d_in_2_a(array_3_io_d_in_2_a),
    .io_d_in_2_valid_a(array_3_io_d_in_2_valid_a),
    .io_d_in_2_b(array_3_io_d_in_2_b),
    .io_d_in_3_a(array_3_io_d_in_3_a),
    .io_d_in_3_valid_a(array_3_io_d_in_3_valid_a),
    .io_d_in_3_b(array_3_io_d_in_3_b),
    .io_d_in_4_a(array_3_io_d_in_4_a),
    .io_d_in_4_valid_a(array_3_io_d_in_4_valid_a),
    .io_d_in_4_b(array_3_io_d_in_4_b),
    .io_d_in_5_a(array_3_io_d_in_5_a),
    .io_d_in_5_valid_a(array_3_io_d_in_5_valid_a),
    .io_d_in_5_b(array_3_io_d_in_5_b),
    .io_d_in_6_a(array_3_io_d_in_6_a),
    .io_d_in_6_valid_a(array_3_io_d_in_6_valid_a),
    .io_d_in_6_b(array_3_io_d_in_6_b),
    .io_d_in_7_a(array_3_io_d_in_7_a),
    .io_d_in_7_valid_a(array_3_io_d_in_7_valid_a),
    .io_d_in_7_b(array_3_io_d_in_7_b),
    .io_d_in_8_a(array_3_io_d_in_8_a),
    .io_d_in_8_valid_a(array_3_io_d_in_8_valid_a),
    .io_d_in_8_b(array_3_io_d_in_8_b),
    .io_d_in_9_a(array_3_io_d_in_9_a),
    .io_d_in_9_valid_a(array_3_io_d_in_9_valid_a),
    .io_d_in_9_b(array_3_io_d_in_9_b),
    .io_d_in_10_a(array_3_io_d_in_10_a),
    .io_d_in_10_valid_a(array_3_io_d_in_10_valid_a),
    .io_d_in_10_b(array_3_io_d_in_10_b),
    .io_d_in_11_a(array_3_io_d_in_11_a),
    .io_d_in_11_valid_a(array_3_io_d_in_11_valid_a),
    .io_d_in_11_b(array_3_io_d_in_11_b),
    .io_d_in_12_a(array_3_io_d_in_12_a),
    .io_d_in_12_valid_a(array_3_io_d_in_12_valid_a),
    .io_d_in_12_b(array_3_io_d_in_12_b),
    .io_d_in_13_a(array_3_io_d_in_13_a),
    .io_d_in_13_valid_a(array_3_io_d_in_13_valid_a),
    .io_d_in_13_b(array_3_io_d_in_13_b),
    .io_d_in_14_a(array_3_io_d_in_14_a),
    .io_d_in_14_valid_a(array_3_io_d_in_14_valid_a),
    .io_d_in_14_b(array_3_io_d_in_14_b),
    .io_d_in_15_a(array_3_io_d_in_15_a),
    .io_d_in_15_valid_a(array_3_io_d_in_15_valid_a),
    .io_d_in_15_b(array_3_io_d_in_15_b),
    .io_d_in_16_a(array_3_io_d_in_16_a),
    .io_d_in_16_valid_a(array_3_io_d_in_16_valid_a),
    .io_d_in_16_b(array_3_io_d_in_16_b),
    .io_d_in_17_a(array_3_io_d_in_17_a),
    .io_d_in_17_valid_a(array_3_io_d_in_17_valid_a),
    .io_d_in_17_b(array_3_io_d_in_17_b),
    .io_d_in_18_a(array_3_io_d_in_18_a),
    .io_d_in_18_valid_a(array_3_io_d_in_18_valid_a),
    .io_d_in_18_b(array_3_io_d_in_18_b),
    .io_d_in_19_a(array_3_io_d_in_19_a),
    .io_d_in_19_valid_a(array_3_io_d_in_19_valid_a),
    .io_d_in_19_b(array_3_io_d_in_19_b),
    .io_d_in_20_a(array_3_io_d_in_20_a),
    .io_d_in_20_valid_a(array_3_io_d_in_20_valid_a),
    .io_d_in_20_b(array_3_io_d_in_20_b),
    .io_d_in_21_a(array_3_io_d_in_21_a),
    .io_d_in_21_valid_a(array_3_io_d_in_21_valid_a),
    .io_d_in_21_b(array_3_io_d_in_21_b),
    .io_d_in_22_a(array_3_io_d_in_22_a),
    .io_d_in_22_valid_a(array_3_io_d_in_22_valid_a),
    .io_d_in_22_b(array_3_io_d_in_22_b),
    .io_d_in_23_a(array_3_io_d_in_23_a),
    .io_d_in_23_valid_a(array_3_io_d_in_23_valid_a),
    .io_d_in_23_b(array_3_io_d_in_23_b),
    .io_d_in_24_a(array_3_io_d_in_24_a),
    .io_d_in_24_valid_a(array_3_io_d_in_24_valid_a),
    .io_d_in_24_b(array_3_io_d_in_24_b),
    .io_d_in_25_a(array_3_io_d_in_25_a),
    .io_d_in_25_valid_a(array_3_io_d_in_25_valid_a),
    .io_d_in_25_b(array_3_io_d_in_25_b),
    .io_d_in_26_a(array_3_io_d_in_26_a),
    .io_d_in_26_valid_a(array_3_io_d_in_26_valid_a),
    .io_d_in_26_b(array_3_io_d_in_26_b),
    .io_d_in_27_a(array_3_io_d_in_27_a),
    .io_d_in_27_valid_a(array_3_io_d_in_27_valid_a),
    .io_d_in_27_b(array_3_io_d_in_27_b),
    .io_d_in_28_a(array_3_io_d_in_28_a),
    .io_d_in_28_valid_a(array_3_io_d_in_28_valid_a),
    .io_d_in_28_b(array_3_io_d_in_28_b),
    .io_d_in_29_a(array_3_io_d_in_29_a),
    .io_d_in_29_valid_a(array_3_io_d_in_29_valid_a),
    .io_d_in_29_b(array_3_io_d_in_29_b),
    .io_d_in_30_a(array_3_io_d_in_30_a),
    .io_d_in_30_valid_a(array_3_io_d_in_30_valid_a),
    .io_d_in_30_b(array_3_io_d_in_30_b),
    .io_d_in_31_a(array_3_io_d_in_31_a),
    .io_d_in_31_valid_a(array_3_io_d_in_31_valid_a),
    .io_d_in_31_b(array_3_io_d_in_31_b),
    .io_d_out_0_a(array_3_io_d_out_0_a),
    .io_d_out_0_valid_a(array_3_io_d_out_0_valid_a),
    .io_d_out_0_b(array_3_io_d_out_0_b),
    .io_d_out_0_valid_b(array_3_io_d_out_0_valid_b),
    .io_d_out_1_a(array_3_io_d_out_1_a),
    .io_d_out_1_valid_a(array_3_io_d_out_1_valid_a),
    .io_d_out_1_b(array_3_io_d_out_1_b),
    .io_d_out_1_valid_b(array_3_io_d_out_1_valid_b),
    .io_d_out_2_a(array_3_io_d_out_2_a),
    .io_d_out_2_valid_a(array_3_io_d_out_2_valid_a),
    .io_d_out_2_b(array_3_io_d_out_2_b),
    .io_d_out_2_valid_b(array_3_io_d_out_2_valid_b),
    .io_d_out_3_a(array_3_io_d_out_3_a),
    .io_d_out_3_valid_a(array_3_io_d_out_3_valid_a),
    .io_d_out_3_b(array_3_io_d_out_3_b),
    .io_d_out_3_valid_b(array_3_io_d_out_3_valid_b),
    .io_d_out_4_a(array_3_io_d_out_4_a),
    .io_d_out_4_valid_a(array_3_io_d_out_4_valid_a),
    .io_d_out_4_b(array_3_io_d_out_4_b),
    .io_d_out_4_valid_b(array_3_io_d_out_4_valid_b),
    .io_d_out_5_a(array_3_io_d_out_5_a),
    .io_d_out_5_valid_a(array_3_io_d_out_5_valid_a),
    .io_d_out_5_b(array_3_io_d_out_5_b),
    .io_d_out_5_valid_b(array_3_io_d_out_5_valid_b),
    .io_d_out_6_a(array_3_io_d_out_6_a),
    .io_d_out_6_valid_a(array_3_io_d_out_6_valid_a),
    .io_d_out_6_b(array_3_io_d_out_6_b),
    .io_d_out_6_valid_b(array_3_io_d_out_6_valid_b),
    .io_d_out_7_a(array_3_io_d_out_7_a),
    .io_d_out_7_valid_a(array_3_io_d_out_7_valid_a),
    .io_d_out_7_b(array_3_io_d_out_7_b),
    .io_d_out_7_valid_b(array_3_io_d_out_7_valid_b),
    .io_d_out_8_a(array_3_io_d_out_8_a),
    .io_d_out_8_valid_a(array_3_io_d_out_8_valid_a),
    .io_d_out_8_b(array_3_io_d_out_8_b),
    .io_d_out_8_valid_b(array_3_io_d_out_8_valid_b),
    .io_d_out_9_a(array_3_io_d_out_9_a),
    .io_d_out_9_valid_a(array_3_io_d_out_9_valid_a),
    .io_d_out_9_b(array_3_io_d_out_9_b),
    .io_d_out_9_valid_b(array_3_io_d_out_9_valid_b),
    .io_d_out_10_a(array_3_io_d_out_10_a),
    .io_d_out_10_valid_a(array_3_io_d_out_10_valid_a),
    .io_d_out_10_b(array_3_io_d_out_10_b),
    .io_d_out_10_valid_b(array_3_io_d_out_10_valid_b),
    .io_d_out_11_a(array_3_io_d_out_11_a),
    .io_d_out_11_valid_a(array_3_io_d_out_11_valid_a),
    .io_d_out_11_b(array_3_io_d_out_11_b),
    .io_d_out_11_valid_b(array_3_io_d_out_11_valid_b),
    .io_d_out_12_a(array_3_io_d_out_12_a),
    .io_d_out_12_valid_a(array_3_io_d_out_12_valid_a),
    .io_d_out_12_b(array_3_io_d_out_12_b),
    .io_d_out_12_valid_b(array_3_io_d_out_12_valid_b),
    .io_d_out_13_a(array_3_io_d_out_13_a),
    .io_d_out_13_valid_a(array_3_io_d_out_13_valid_a),
    .io_d_out_13_b(array_3_io_d_out_13_b),
    .io_d_out_13_valid_b(array_3_io_d_out_13_valid_b),
    .io_d_out_14_a(array_3_io_d_out_14_a),
    .io_d_out_14_valid_a(array_3_io_d_out_14_valid_a),
    .io_d_out_14_b(array_3_io_d_out_14_b),
    .io_d_out_14_valid_b(array_3_io_d_out_14_valid_b),
    .io_d_out_15_a(array_3_io_d_out_15_a),
    .io_d_out_15_valid_a(array_3_io_d_out_15_valid_a),
    .io_d_out_15_b(array_3_io_d_out_15_b),
    .io_d_out_15_valid_b(array_3_io_d_out_15_valid_b),
    .io_d_out_16_a(array_3_io_d_out_16_a),
    .io_d_out_16_valid_a(array_3_io_d_out_16_valid_a),
    .io_d_out_16_b(array_3_io_d_out_16_b),
    .io_d_out_16_valid_b(array_3_io_d_out_16_valid_b),
    .io_d_out_17_a(array_3_io_d_out_17_a),
    .io_d_out_17_valid_a(array_3_io_d_out_17_valid_a),
    .io_d_out_17_b(array_3_io_d_out_17_b),
    .io_d_out_17_valid_b(array_3_io_d_out_17_valid_b),
    .io_d_out_18_a(array_3_io_d_out_18_a),
    .io_d_out_18_valid_a(array_3_io_d_out_18_valid_a),
    .io_d_out_18_b(array_3_io_d_out_18_b),
    .io_d_out_18_valid_b(array_3_io_d_out_18_valid_b),
    .io_d_out_19_a(array_3_io_d_out_19_a),
    .io_d_out_19_valid_a(array_3_io_d_out_19_valid_a),
    .io_d_out_19_b(array_3_io_d_out_19_b),
    .io_d_out_19_valid_b(array_3_io_d_out_19_valid_b),
    .io_d_out_20_a(array_3_io_d_out_20_a),
    .io_d_out_20_valid_a(array_3_io_d_out_20_valid_a),
    .io_d_out_20_b(array_3_io_d_out_20_b),
    .io_d_out_20_valid_b(array_3_io_d_out_20_valid_b),
    .io_d_out_21_a(array_3_io_d_out_21_a),
    .io_d_out_21_valid_a(array_3_io_d_out_21_valid_a),
    .io_d_out_21_b(array_3_io_d_out_21_b),
    .io_d_out_21_valid_b(array_3_io_d_out_21_valid_b),
    .io_d_out_22_a(array_3_io_d_out_22_a),
    .io_d_out_22_valid_a(array_3_io_d_out_22_valid_a),
    .io_d_out_22_b(array_3_io_d_out_22_b),
    .io_d_out_22_valid_b(array_3_io_d_out_22_valid_b),
    .io_d_out_23_a(array_3_io_d_out_23_a),
    .io_d_out_23_valid_a(array_3_io_d_out_23_valid_a),
    .io_d_out_23_b(array_3_io_d_out_23_b),
    .io_d_out_23_valid_b(array_3_io_d_out_23_valid_b),
    .io_d_out_24_a(array_3_io_d_out_24_a),
    .io_d_out_24_valid_a(array_3_io_d_out_24_valid_a),
    .io_d_out_24_b(array_3_io_d_out_24_b),
    .io_d_out_24_valid_b(array_3_io_d_out_24_valid_b),
    .io_d_out_25_a(array_3_io_d_out_25_a),
    .io_d_out_25_valid_a(array_3_io_d_out_25_valid_a),
    .io_d_out_25_b(array_3_io_d_out_25_b),
    .io_d_out_25_valid_b(array_3_io_d_out_25_valid_b),
    .io_d_out_26_a(array_3_io_d_out_26_a),
    .io_d_out_26_valid_a(array_3_io_d_out_26_valid_a),
    .io_d_out_26_b(array_3_io_d_out_26_b),
    .io_d_out_26_valid_b(array_3_io_d_out_26_valid_b),
    .io_d_out_27_a(array_3_io_d_out_27_a),
    .io_d_out_27_valid_a(array_3_io_d_out_27_valid_a),
    .io_d_out_27_b(array_3_io_d_out_27_b),
    .io_d_out_27_valid_b(array_3_io_d_out_27_valid_b),
    .io_d_out_28_a(array_3_io_d_out_28_a),
    .io_d_out_28_valid_a(array_3_io_d_out_28_valid_a),
    .io_d_out_28_b(array_3_io_d_out_28_b),
    .io_d_out_28_valid_b(array_3_io_d_out_28_valid_b),
    .io_d_out_29_a(array_3_io_d_out_29_a),
    .io_d_out_29_valid_a(array_3_io_d_out_29_valid_a),
    .io_d_out_29_b(array_3_io_d_out_29_b),
    .io_d_out_29_valid_b(array_3_io_d_out_29_valid_b),
    .io_d_out_30_a(array_3_io_d_out_30_a),
    .io_d_out_30_valid_a(array_3_io_d_out_30_valid_a),
    .io_d_out_30_b(array_3_io_d_out_30_b),
    .io_d_out_30_valid_b(array_3_io_d_out_30_valid_b),
    .io_d_out_31_a(array_3_io_d_out_31_a),
    .io_d_out_31_valid_a(array_3_io_d_out_31_valid_a),
    .io_d_out_31_b(array_3_io_d_out_31_b),
    .io_d_out_31_valid_b(array_3_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_3_io_wr_en_mem1),
    .io_wr_en_mem2(array_3_io_wr_en_mem2),
    .io_wr_en_mem3(array_3_io_wr_en_mem3),
    .io_wr_en_mem4(array_3_io_wr_en_mem4),
    .io_wr_en_mem5(array_3_io_wr_en_mem5),
    .io_wr_en_mem6(array_3_io_wr_en_mem6),
    .io_wr_instr_mem1(array_3_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_3_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_3_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_3_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_3_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_3_io_wr_instr_mem6),
    .io_PC1_in(array_3_io_PC1_in),
    .io_PC6_out(array_3_io_PC6_out),
    .io_Addr_in(array_3_io_Addr_in),
    .io_Addr_out(array_3_io_Addr_out),
    .io_Tag_in_Tag(array_3_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_3_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_3_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_3_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_4 ( // @[Array.scala 41:54]
    .clock(array_4_clock),
    .reset(array_4_reset),
    .io_d_in_0_a(array_4_io_d_in_0_a),
    .io_d_in_0_valid_a(array_4_io_d_in_0_valid_a),
    .io_d_in_0_b(array_4_io_d_in_0_b),
    .io_d_in_1_a(array_4_io_d_in_1_a),
    .io_d_in_1_valid_a(array_4_io_d_in_1_valid_a),
    .io_d_in_1_b(array_4_io_d_in_1_b),
    .io_d_in_2_a(array_4_io_d_in_2_a),
    .io_d_in_2_valid_a(array_4_io_d_in_2_valid_a),
    .io_d_in_2_b(array_4_io_d_in_2_b),
    .io_d_in_3_a(array_4_io_d_in_3_a),
    .io_d_in_3_valid_a(array_4_io_d_in_3_valid_a),
    .io_d_in_3_b(array_4_io_d_in_3_b),
    .io_d_in_4_a(array_4_io_d_in_4_a),
    .io_d_in_4_valid_a(array_4_io_d_in_4_valid_a),
    .io_d_in_4_b(array_4_io_d_in_4_b),
    .io_d_in_5_a(array_4_io_d_in_5_a),
    .io_d_in_5_valid_a(array_4_io_d_in_5_valid_a),
    .io_d_in_5_b(array_4_io_d_in_5_b),
    .io_d_in_6_a(array_4_io_d_in_6_a),
    .io_d_in_6_valid_a(array_4_io_d_in_6_valid_a),
    .io_d_in_6_b(array_4_io_d_in_6_b),
    .io_d_in_7_a(array_4_io_d_in_7_a),
    .io_d_in_7_valid_a(array_4_io_d_in_7_valid_a),
    .io_d_in_7_b(array_4_io_d_in_7_b),
    .io_d_in_8_a(array_4_io_d_in_8_a),
    .io_d_in_8_valid_a(array_4_io_d_in_8_valid_a),
    .io_d_in_8_b(array_4_io_d_in_8_b),
    .io_d_in_9_a(array_4_io_d_in_9_a),
    .io_d_in_9_valid_a(array_4_io_d_in_9_valid_a),
    .io_d_in_9_b(array_4_io_d_in_9_b),
    .io_d_in_10_a(array_4_io_d_in_10_a),
    .io_d_in_10_valid_a(array_4_io_d_in_10_valid_a),
    .io_d_in_10_b(array_4_io_d_in_10_b),
    .io_d_in_11_a(array_4_io_d_in_11_a),
    .io_d_in_11_valid_a(array_4_io_d_in_11_valid_a),
    .io_d_in_11_b(array_4_io_d_in_11_b),
    .io_d_in_12_a(array_4_io_d_in_12_a),
    .io_d_in_12_valid_a(array_4_io_d_in_12_valid_a),
    .io_d_in_12_b(array_4_io_d_in_12_b),
    .io_d_in_13_a(array_4_io_d_in_13_a),
    .io_d_in_13_valid_a(array_4_io_d_in_13_valid_a),
    .io_d_in_13_b(array_4_io_d_in_13_b),
    .io_d_in_14_a(array_4_io_d_in_14_a),
    .io_d_in_14_valid_a(array_4_io_d_in_14_valid_a),
    .io_d_in_14_b(array_4_io_d_in_14_b),
    .io_d_in_15_a(array_4_io_d_in_15_a),
    .io_d_in_15_valid_a(array_4_io_d_in_15_valid_a),
    .io_d_in_15_b(array_4_io_d_in_15_b),
    .io_d_in_16_a(array_4_io_d_in_16_a),
    .io_d_in_16_valid_a(array_4_io_d_in_16_valid_a),
    .io_d_in_16_b(array_4_io_d_in_16_b),
    .io_d_in_17_a(array_4_io_d_in_17_a),
    .io_d_in_17_valid_a(array_4_io_d_in_17_valid_a),
    .io_d_in_17_b(array_4_io_d_in_17_b),
    .io_d_in_18_a(array_4_io_d_in_18_a),
    .io_d_in_18_valid_a(array_4_io_d_in_18_valid_a),
    .io_d_in_18_b(array_4_io_d_in_18_b),
    .io_d_in_19_a(array_4_io_d_in_19_a),
    .io_d_in_19_valid_a(array_4_io_d_in_19_valid_a),
    .io_d_in_19_b(array_4_io_d_in_19_b),
    .io_d_in_20_a(array_4_io_d_in_20_a),
    .io_d_in_20_valid_a(array_4_io_d_in_20_valid_a),
    .io_d_in_20_b(array_4_io_d_in_20_b),
    .io_d_in_21_a(array_4_io_d_in_21_a),
    .io_d_in_21_valid_a(array_4_io_d_in_21_valid_a),
    .io_d_in_21_b(array_4_io_d_in_21_b),
    .io_d_in_22_a(array_4_io_d_in_22_a),
    .io_d_in_22_valid_a(array_4_io_d_in_22_valid_a),
    .io_d_in_22_b(array_4_io_d_in_22_b),
    .io_d_in_23_a(array_4_io_d_in_23_a),
    .io_d_in_23_valid_a(array_4_io_d_in_23_valid_a),
    .io_d_in_23_b(array_4_io_d_in_23_b),
    .io_d_in_24_a(array_4_io_d_in_24_a),
    .io_d_in_24_valid_a(array_4_io_d_in_24_valid_a),
    .io_d_in_24_b(array_4_io_d_in_24_b),
    .io_d_in_25_a(array_4_io_d_in_25_a),
    .io_d_in_25_valid_a(array_4_io_d_in_25_valid_a),
    .io_d_in_25_b(array_4_io_d_in_25_b),
    .io_d_in_26_a(array_4_io_d_in_26_a),
    .io_d_in_26_valid_a(array_4_io_d_in_26_valid_a),
    .io_d_in_26_b(array_4_io_d_in_26_b),
    .io_d_in_27_a(array_4_io_d_in_27_a),
    .io_d_in_27_valid_a(array_4_io_d_in_27_valid_a),
    .io_d_in_27_b(array_4_io_d_in_27_b),
    .io_d_in_28_a(array_4_io_d_in_28_a),
    .io_d_in_28_valid_a(array_4_io_d_in_28_valid_a),
    .io_d_in_28_b(array_4_io_d_in_28_b),
    .io_d_in_29_a(array_4_io_d_in_29_a),
    .io_d_in_29_valid_a(array_4_io_d_in_29_valid_a),
    .io_d_in_29_b(array_4_io_d_in_29_b),
    .io_d_in_30_a(array_4_io_d_in_30_a),
    .io_d_in_30_valid_a(array_4_io_d_in_30_valid_a),
    .io_d_in_30_b(array_4_io_d_in_30_b),
    .io_d_in_31_a(array_4_io_d_in_31_a),
    .io_d_in_31_valid_a(array_4_io_d_in_31_valid_a),
    .io_d_in_31_b(array_4_io_d_in_31_b),
    .io_d_out_0_a(array_4_io_d_out_0_a),
    .io_d_out_0_valid_a(array_4_io_d_out_0_valid_a),
    .io_d_out_0_b(array_4_io_d_out_0_b),
    .io_d_out_0_valid_b(array_4_io_d_out_0_valid_b),
    .io_d_out_1_a(array_4_io_d_out_1_a),
    .io_d_out_1_valid_a(array_4_io_d_out_1_valid_a),
    .io_d_out_1_b(array_4_io_d_out_1_b),
    .io_d_out_1_valid_b(array_4_io_d_out_1_valid_b),
    .io_d_out_2_a(array_4_io_d_out_2_a),
    .io_d_out_2_valid_a(array_4_io_d_out_2_valid_a),
    .io_d_out_2_b(array_4_io_d_out_2_b),
    .io_d_out_2_valid_b(array_4_io_d_out_2_valid_b),
    .io_d_out_3_a(array_4_io_d_out_3_a),
    .io_d_out_3_valid_a(array_4_io_d_out_3_valid_a),
    .io_d_out_3_b(array_4_io_d_out_3_b),
    .io_d_out_3_valid_b(array_4_io_d_out_3_valid_b),
    .io_d_out_4_a(array_4_io_d_out_4_a),
    .io_d_out_4_valid_a(array_4_io_d_out_4_valid_a),
    .io_d_out_4_b(array_4_io_d_out_4_b),
    .io_d_out_4_valid_b(array_4_io_d_out_4_valid_b),
    .io_d_out_5_a(array_4_io_d_out_5_a),
    .io_d_out_5_valid_a(array_4_io_d_out_5_valid_a),
    .io_d_out_5_b(array_4_io_d_out_5_b),
    .io_d_out_5_valid_b(array_4_io_d_out_5_valid_b),
    .io_d_out_6_a(array_4_io_d_out_6_a),
    .io_d_out_6_valid_a(array_4_io_d_out_6_valid_a),
    .io_d_out_6_b(array_4_io_d_out_6_b),
    .io_d_out_6_valid_b(array_4_io_d_out_6_valid_b),
    .io_d_out_7_a(array_4_io_d_out_7_a),
    .io_d_out_7_valid_a(array_4_io_d_out_7_valid_a),
    .io_d_out_7_b(array_4_io_d_out_7_b),
    .io_d_out_7_valid_b(array_4_io_d_out_7_valid_b),
    .io_d_out_8_a(array_4_io_d_out_8_a),
    .io_d_out_8_valid_a(array_4_io_d_out_8_valid_a),
    .io_d_out_8_b(array_4_io_d_out_8_b),
    .io_d_out_8_valid_b(array_4_io_d_out_8_valid_b),
    .io_d_out_9_a(array_4_io_d_out_9_a),
    .io_d_out_9_valid_a(array_4_io_d_out_9_valid_a),
    .io_d_out_9_b(array_4_io_d_out_9_b),
    .io_d_out_9_valid_b(array_4_io_d_out_9_valid_b),
    .io_d_out_10_a(array_4_io_d_out_10_a),
    .io_d_out_10_valid_a(array_4_io_d_out_10_valid_a),
    .io_d_out_10_b(array_4_io_d_out_10_b),
    .io_d_out_10_valid_b(array_4_io_d_out_10_valid_b),
    .io_d_out_11_a(array_4_io_d_out_11_a),
    .io_d_out_11_valid_a(array_4_io_d_out_11_valid_a),
    .io_d_out_11_b(array_4_io_d_out_11_b),
    .io_d_out_11_valid_b(array_4_io_d_out_11_valid_b),
    .io_d_out_12_a(array_4_io_d_out_12_a),
    .io_d_out_12_valid_a(array_4_io_d_out_12_valid_a),
    .io_d_out_12_b(array_4_io_d_out_12_b),
    .io_d_out_12_valid_b(array_4_io_d_out_12_valid_b),
    .io_d_out_13_a(array_4_io_d_out_13_a),
    .io_d_out_13_valid_a(array_4_io_d_out_13_valid_a),
    .io_d_out_13_b(array_4_io_d_out_13_b),
    .io_d_out_13_valid_b(array_4_io_d_out_13_valid_b),
    .io_d_out_14_a(array_4_io_d_out_14_a),
    .io_d_out_14_valid_a(array_4_io_d_out_14_valid_a),
    .io_d_out_14_b(array_4_io_d_out_14_b),
    .io_d_out_14_valid_b(array_4_io_d_out_14_valid_b),
    .io_d_out_15_a(array_4_io_d_out_15_a),
    .io_d_out_15_valid_a(array_4_io_d_out_15_valid_a),
    .io_d_out_15_b(array_4_io_d_out_15_b),
    .io_d_out_15_valid_b(array_4_io_d_out_15_valid_b),
    .io_d_out_16_a(array_4_io_d_out_16_a),
    .io_d_out_16_valid_a(array_4_io_d_out_16_valid_a),
    .io_d_out_16_b(array_4_io_d_out_16_b),
    .io_d_out_16_valid_b(array_4_io_d_out_16_valid_b),
    .io_d_out_17_a(array_4_io_d_out_17_a),
    .io_d_out_17_valid_a(array_4_io_d_out_17_valid_a),
    .io_d_out_17_b(array_4_io_d_out_17_b),
    .io_d_out_17_valid_b(array_4_io_d_out_17_valid_b),
    .io_d_out_18_a(array_4_io_d_out_18_a),
    .io_d_out_18_valid_a(array_4_io_d_out_18_valid_a),
    .io_d_out_18_b(array_4_io_d_out_18_b),
    .io_d_out_18_valid_b(array_4_io_d_out_18_valid_b),
    .io_d_out_19_a(array_4_io_d_out_19_a),
    .io_d_out_19_valid_a(array_4_io_d_out_19_valid_a),
    .io_d_out_19_b(array_4_io_d_out_19_b),
    .io_d_out_19_valid_b(array_4_io_d_out_19_valid_b),
    .io_d_out_20_a(array_4_io_d_out_20_a),
    .io_d_out_20_valid_a(array_4_io_d_out_20_valid_a),
    .io_d_out_20_b(array_4_io_d_out_20_b),
    .io_d_out_20_valid_b(array_4_io_d_out_20_valid_b),
    .io_d_out_21_a(array_4_io_d_out_21_a),
    .io_d_out_21_valid_a(array_4_io_d_out_21_valid_a),
    .io_d_out_21_b(array_4_io_d_out_21_b),
    .io_d_out_21_valid_b(array_4_io_d_out_21_valid_b),
    .io_d_out_22_a(array_4_io_d_out_22_a),
    .io_d_out_22_valid_a(array_4_io_d_out_22_valid_a),
    .io_d_out_22_b(array_4_io_d_out_22_b),
    .io_d_out_22_valid_b(array_4_io_d_out_22_valid_b),
    .io_d_out_23_a(array_4_io_d_out_23_a),
    .io_d_out_23_valid_a(array_4_io_d_out_23_valid_a),
    .io_d_out_23_b(array_4_io_d_out_23_b),
    .io_d_out_23_valid_b(array_4_io_d_out_23_valid_b),
    .io_d_out_24_a(array_4_io_d_out_24_a),
    .io_d_out_24_valid_a(array_4_io_d_out_24_valid_a),
    .io_d_out_24_b(array_4_io_d_out_24_b),
    .io_d_out_24_valid_b(array_4_io_d_out_24_valid_b),
    .io_d_out_25_a(array_4_io_d_out_25_a),
    .io_d_out_25_valid_a(array_4_io_d_out_25_valid_a),
    .io_d_out_25_b(array_4_io_d_out_25_b),
    .io_d_out_25_valid_b(array_4_io_d_out_25_valid_b),
    .io_d_out_26_a(array_4_io_d_out_26_a),
    .io_d_out_26_valid_a(array_4_io_d_out_26_valid_a),
    .io_d_out_26_b(array_4_io_d_out_26_b),
    .io_d_out_26_valid_b(array_4_io_d_out_26_valid_b),
    .io_d_out_27_a(array_4_io_d_out_27_a),
    .io_d_out_27_valid_a(array_4_io_d_out_27_valid_a),
    .io_d_out_27_b(array_4_io_d_out_27_b),
    .io_d_out_27_valid_b(array_4_io_d_out_27_valid_b),
    .io_d_out_28_a(array_4_io_d_out_28_a),
    .io_d_out_28_valid_a(array_4_io_d_out_28_valid_a),
    .io_d_out_28_b(array_4_io_d_out_28_b),
    .io_d_out_28_valid_b(array_4_io_d_out_28_valid_b),
    .io_d_out_29_a(array_4_io_d_out_29_a),
    .io_d_out_29_valid_a(array_4_io_d_out_29_valid_a),
    .io_d_out_29_b(array_4_io_d_out_29_b),
    .io_d_out_29_valid_b(array_4_io_d_out_29_valid_b),
    .io_d_out_30_a(array_4_io_d_out_30_a),
    .io_d_out_30_valid_a(array_4_io_d_out_30_valid_a),
    .io_d_out_30_b(array_4_io_d_out_30_b),
    .io_d_out_30_valid_b(array_4_io_d_out_30_valid_b),
    .io_d_out_31_a(array_4_io_d_out_31_a),
    .io_d_out_31_valid_a(array_4_io_d_out_31_valid_a),
    .io_d_out_31_b(array_4_io_d_out_31_b),
    .io_d_out_31_valid_b(array_4_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_4_io_wr_en_mem1),
    .io_wr_en_mem2(array_4_io_wr_en_mem2),
    .io_wr_en_mem3(array_4_io_wr_en_mem3),
    .io_wr_en_mem4(array_4_io_wr_en_mem4),
    .io_wr_en_mem5(array_4_io_wr_en_mem5),
    .io_wr_en_mem6(array_4_io_wr_en_mem6),
    .io_wr_instr_mem1(array_4_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_4_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_4_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_4_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_4_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_4_io_wr_instr_mem6),
    .io_PC1_in(array_4_io_PC1_in),
    .io_PC6_out(array_4_io_PC6_out),
    .io_Addr_in(array_4_io_Addr_in),
    .io_Addr_out(array_4_io_Addr_out),
    .io_Tag_in_Tag(array_4_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_4_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_4_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_4_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_5 ( // @[Array.scala 41:54]
    .clock(array_5_clock),
    .reset(array_5_reset),
    .io_d_in_0_a(array_5_io_d_in_0_a),
    .io_d_in_0_valid_a(array_5_io_d_in_0_valid_a),
    .io_d_in_0_b(array_5_io_d_in_0_b),
    .io_d_in_1_a(array_5_io_d_in_1_a),
    .io_d_in_1_valid_a(array_5_io_d_in_1_valid_a),
    .io_d_in_1_b(array_5_io_d_in_1_b),
    .io_d_in_2_a(array_5_io_d_in_2_a),
    .io_d_in_2_valid_a(array_5_io_d_in_2_valid_a),
    .io_d_in_2_b(array_5_io_d_in_2_b),
    .io_d_in_3_a(array_5_io_d_in_3_a),
    .io_d_in_3_valid_a(array_5_io_d_in_3_valid_a),
    .io_d_in_3_b(array_5_io_d_in_3_b),
    .io_d_in_4_a(array_5_io_d_in_4_a),
    .io_d_in_4_valid_a(array_5_io_d_in_4_valid_a),
    .io_d_in_4_b(array_5_io_d_in_4_b),
    .io_d_in_5_a(array_5_io_d_in_5_a),
    .io_d_in_5_valid_a(array_5_io_d_in_5_valid_a),
    .io_d_in_5_b(array_5_io_d_in_5_b),
    .io_d_in_6_a(array_5_io_d_in_6_a),
    .io_d_in_6_valid_a(array_5_io_d_in_6_valid_a),
    .io_d_in_6_b(array_5_io_d_in_6_b),
    .io_d_in_7_a(array_5_io_d_in_7_a),
    .io_d_in_7_valid_a(array_5_io_d_in_7_valid_a),
    .io_d_in_7_b(array_5_io_d_in_7_b),
    .io_d_in_8_a(array_5_io_d_in_8_a),
    .io_d_in_8_valid_a(array_5_io_d_in_8_valid_a),
    .io_d_in_8_b(array_5_io_d_in_8_b),
    .io_d_in_9_a(array_5_io_d_in_9_a),
    .io_d_in_9_valid_a(array_5_io_d_in_9_valid_a),
    .io_d_in_9_b(array_5_io_d_in_9_b),
    .io_d_in_10_a(array_5_io_d_in_10_a),
    .io_d_in_10_valid_a(array_5_io_d_in_10_valid_a),
    .io_d_in_10_b(array_5_io_d_in_10_b),
    .io_d_in_11_a(array_5_io_d_in_11_a),
    .io_d_in_11_valid_a(array_5_io_d_in_11_valid_a),
    .io_d_in_11_b(array_5_io_d_in_11_b),
    .io_d_in_12_a(array_5_io_d_in_12_a),
    .io_d_in_12_valid_a(array_5_io_d_in_12_valid_a),
    .io_d_in_12_b(array_5_io_d_in_12_b),
    .io_d_in_13_a(array_5_io_d_in_13_a),
    .io_d_in_13_valid_a(array_5_io_d_in_13_valid_a),
    .io_d_in_13_b(array_5_io_d_in_13_b),
    .io_d_in_14_a(array_5_io_d_in_14_a),
    .io_d_in_14_valid_a(array_5_io_d_in_14_valid_a),
    .io_d_in_14_b(array_5_io_d_in_14_b),
    .io_d_in_15_a(array_5_io_d_in_15_a),
    .io_d_in_15_valid_a(array_5_io_d_in_15_valid_a),
    .io_d_in_15_b(array_5_io_d_in_15_b),
    .io_d_in_16_a(array_5_io_d_in_16_a),
    .io_d_in_16_valid_a(array_5_io_d_in_16_valid_a),
    .io_d_in_16_b(array_5_io_d_in_16_b),
    .io_d_in_17_a(array_5_io_d_in_17_a),
    .io_d_in_17_valid_a(array_5_io_d_in_17_valid_a),
    .io_d_in_17_b(array_5_io_d_in_17_b),
    .io_d_in_18_a(array_5_io_d_in_18_a),
    .io_d_in_18_valid_a(array_5_io_d_in_18_valid_a),
    .io_d_in_18_b(array_5_io_d_in_18_b),
    .io_d_in_19_a(array_5_io_d_in_19_a),
    .io_d_in_19_valid_a(array_5_io_d_in_19_valid_a),
    .io_d_in_19_b(array_5_io_d_in_19_b),
    .io_d_in_20_a(array_5_io_d_in_20_a),
    .io_d_in_20_valid_a(array_5_io_d_in_20_valid_a),
    .io_d_in_20_b(array_5_io_d_in_20_b),
    .io_d_in_21_a(array_5_io_d_in_21_a),
    .io_d_in_21_valid_a(array_5_io_d_in_21_valid_a),
    .io_d_in_21_b(array_5_io_d_in_21_b),
    .io_d_in_22_a(array_5_io_d_in_22_a),
    .io_d_in_22_valid_a(array_5_io_d_in_22_valid_a),
    .io_d_in_22_b(array_5_io_d_in_22_b),
    .io_d_in_23_a(array_5_io_d_in_23_a),
    .io_d_in_23_valid_a(array_5_io_d_in_23_valid_a),
    .io_d_in_23_b(array_5_io_d_in_23_b),
    .io_d_in_24_a(array_5_io_d_in_24_a),
    .io_d_in_24_valid_a(array_5_io_d_in_24_valid_a),
    .io_d_in_24_b(array_5_io_d_in_24_b),
    .io_d_in_25_a(array_5_io_d_in_25_a),
    .io_d_in_25_valid_a(array_5_io_d_in_25_valid_a),
    .io_d_in_25_b(array_5_io_d_in_25_b),
    .io_d_in_26_a(array_5_io_d_in_26_a),
    .io_d_in_26_valid_a(array_5_io_d_in_26_valid_a),
    .io_d_in_26_b(array_5_io_d_in_26_b),
    .io_d_in_27_a(array_5_io_d_in_27_a),
    .io_d_in_27_valid_a(array_5_io_d_in_27_valid_a),
    .io_d_in_27_b(array_5_io_d_in_27_b),
    .io_d_in_28_a(array_5_io_d_in_28_a),
    .io_d_in_28_valid_a(array_5_io_d_in_28_valid_a),
    .io_d_in_28_b(array_5_io_d_in_28_b),
    .io_d_in_29_a(array_5_io_d_in_29_a),
    .io_d_in_29_valid_a(array_5_io_d_in_29_valid_a),
    .io_d_in_29_b(array_5_io_d_in_29_b),
    .io_d_in_30_a(array_5_io_d_in_30_a),
    .io_d_in_30_valid_a(array_5_io_d_in_30_valid_a),
    .io_d_in_30_b(array_5_io_d_in_30_b),
    .io_d_in_31_a(array_5_io_d_in_31_a),
    .io_d_in_31_valid_a(array_5_io_d_in_31_valid_a),
    .io_d_in_31_b(array_5_io_d_in_31_b),
    .io_d_out_0_a(array_5_io_d_out_0_a),
    .io_d_out_0_valid_a(array_5_io_d_out_0_valid_a),
    .io_d_out_0_b(array_5_io_d_out_0_b),
    .io_d_out_0_valid_b(array_5_io_d_out_0_valid_b),
    .io_d_out_1_a(array_5_io_d_out_1_a),
    .io_d_out_1_valid_a(array_5_io_d_out_1_valid_a),
    .io_d_out_1_b(array_5_io_d_out_1_b),
    .io_d_out_1_valid_b(array_5_io_d_out_1_valid_b),
    .io_d_out_2_a(array_5_io_d_out_2_a),
    .io_d_out_2_valid_a(array_5_io_d_out_2_valid_a),
    .io_d_out_2_b(array_5_io_d_out_2_b),
    .io_d_out_2_valid_b(array_5_io_d_out_2_valid_b),
    .io_d_out_3_a(array_5_io_d_out_3_a),
    .io_d_out_3_valid_a(array_5_io_d_out_3_valid_a),
    .io_d_out_3_b(array_5_io_d_out_3_b),
    .io_d_out_3_valid_b(array_5_io_d_out_3_valid_b),
    .io_d_out_4_a(array_5_io_d_out_4_a),
    .io_d_out_4_valid_a(array_5_io_d_out_4_valid_a),
    .io_d_out_4_b(array_5_io_d_out_4_b),
    .io_d_out_4_valid_b(array_5_io_d_out_4_valid_b),
    .io_d_out_5_a(array_5_io_d_out_5_a),
    .io_d_out_5_valid_a(array_5_io_d_out_5_valid_a),
    .io_d_out_5_b(array_5_io_d_out_5_b),
    .io_d_out_5_valid_b(array_5_io_d_out_5_valid_b),
    .io_d_out_6_a(array_5_io_d_out_6_a),
    .io_d_out_6_valid_a(array_5_io_d_out_6_valid_a),
    .io_d_out_6_b(array_5_io_d_out_6_b),
    .io_d_out_6_valid_b(array_5_io_d_out_6_valid_b),
    .io_d_out_7_a(array_5_io_d_out_7_a),
    .io_d_out_7_valid_a(array_5_io_d_out_7_valid_a),
    .io_d_out_7_b(array_5_io_d_out_7_b),
    .io_d_out_7_valid_b(array_5_io_d_out_7_valid_b),
    .io_d_out_8_a(array_5_io_d_out_8_a),
    .io_d_out_8_valid_a(array_5_io_d_out_8_valid_a),
    .io_d_out_8_b(array_5_io_d_out_8_b),
    .io_d_out_8_valid_b(array_5_io_d_out_8_valid_b),
    .io_d_out_9_a(array_5_io_d_out_9_a),
    .io_d_out_9_valid_a(array_5_io_d_out_9_valid_a),
    .io_d_out_9_b(array_5_io_d_out_9_b),
    .io_d_out_9_valid_b(array_5_io_d_out_9_valid_b),
    .io_d_out_10_a(array_5_io_d_out_10_a),
    .io_d_out_10_valid_a(array_5_io_d_out_10_valid_a),
    .io_d_out_10_b(array_5_io_d_out_10_b),
    .io_d_out_10_valid_b(array_5_io_d_out_10_valid_b),
    .io_d_out_11_a(array_5_io_d_out_11_a),
    .io_d_out_11_valid_a(array_5_io_d_out_11_valid_a),
    .io_d_out_11_b(array_5_io_d_out_11_b),
    .io_d_out_11_valid_b(array_5_io_d_out_11_valid_b),
    .io_d_out_12_a(array_5_io_d_out_12_a),
    .io_d_out_12_valid_a(array_5_io_d_out_12_valid_a),
    .io_d_out_12_b(array_5_io_d_out_12_b),
    .io_d_out_12_valid_b(array_5_io_d_out_12_valid_b),
    .io_d_out_13_a(array_5_io_d_out_13_a),
    .io_d_out_13_valid_a(array_5_io_d_out_13_valid_a),
    .io_d_out_13_b(array_5_io_d_out_13_b),
    .io_d_out_13_valid_b(array_5_io_d_out_13_valid_b),
    .io_d_out_14_a(array_5_io_d_out_14_a),
    .io_d_out_14_valid_a(array_5_io_d_out_14_valid_a),
    .io_d_out_14_b(array_5_io_d_out_14_b),
    .io_d_out_14_valid_b(array_5_io_d_out_14_valid_b),
    .io_d_out_15_a(array_5_io_d_out_15_a),
    .io_d_out_15_valid_a(array_5_io_d_out_15_valid_a),
    .io_d_out_15_b(array_5_io_d_out_15_b),
    .io_d_out_15_valid_b(array_5_io_d_out_15_valid_b),
    .io_d_out_16_a(array_5_io_d_out_16_a),
    .io_d_out_16_valid_a(array_5_io_d_out_16_valid_a),
    .io_d_out_16_b(array_5_io_d_out_16_b),
    .io_d_out_16_valid_b(array_5_io_d_out_16_valid_b),
    .io_d_out_17_a(array_5_io_d_out_17_a),
    .io_d_out_17_valid_a(array_5_io_d_out_17_valid_a),
    .io_d_out_17_b(array_5_io_d_out_17_b),
    .io_d_out_17_valid_b(array_5_io_d_out_17_valid_b),
    .io_d_out_18_a(array_5_io_d_out_18_a),
    .io_d_out_18_valid_a(array_5_io_d_out_18_valid_a),
    .io_d_out_18_b(array_5_io_d_out_18_b),
    .io_d_out_18_valid_b(array_5_io_d_out_18_valid_b),
    .io_d_out_19_a(array_5_io_d_out_19_a),
    .io_d_out_19_valid_a(array_5_io_d_out_19_valid_a),
    .io_d_out_19_b(array_5_io_d_out_19_b),
    .io_d_out_19_valid_b(array_5_io_d_out_19_valid_b),
    .io_d_out_20_a(array_5_io_d_out_20_a),
    .io_d_out_20_valid_a(array_5_io_d_out_20_valid_a),
    .io_d_out_20_b(array_5_io_d_out_20_b),
    .io_d_out_20_valid_b(array_5_io_d_out_20_valid_b),
    .io_d_out_21_a(array_5_io_d_out_21_a),
    .io_d_out_21_valid_a(array_5_io_d_out_21_valid_a),
    .io_d_out_21_b(array_5_io_d_out_21_b),
    .io_d_out_21_valid_b(array_5_io_d_out_21_valid_b),
    .io_d_out_22_a(array_5_io_d_out_22_a),
    .io_d_out_22_valid_a(array_5_io_d_out_22_valid_a),
    .io_d_out_22_b(array_5_io_d_out_22_b),
    .io_d_out_22_valid_b(array_5_io_d_out_22_valid_b),
    .io_d_out_23_a(array_5_io_d_out_23_a),
    .io_d_out_23_valid_a(array_5_io_d_out_23_valid_a),
    .io_d_out_23_b(array_5_io_d_out_23_b),
    .io_d_out_23_valid_b(array_5_io_d_out_23_valid_b),
    .io_d_out_24_a(array_5_io_d_out_24_a),
    .io_d_out_24_valid_a(array_5_io_d_out_24_valid_a),
    .io_d_out_24_b(array_5_io_d_out_24_b),
    .io_d_out_24_valid_b(array_5_io_d_out_24_valid_b),
    .io_d_out_25_a(array_5_io_d_out_25_a),
    .io_d_out_25_valid_a(array_5_io_d_out_25_valid_a),
    .io_d_out_25_b(array_5_io_d_out_25_b),
    .io_d_out_25_valid_b(array_5_io_d_out_25_valid_b),
    .io_d_out_26_a(array_5_io_d_out_26_a),
    .io_d_out_26_valid_a(array_5_io_d_out_26_valid_a),
    .io_d_out_26_b(array_5_io_d_out_26_b),
    .io_d_out_26_valid_b(array_5_io_d_out_26_valid_b),
    .io_d_out_27_a(array_5_io_d_out_27_a),
    .io_d_out_27_valid_a(array_5_io_d_out_27_valid_a),
    .io_d_out_27_b(array_5_io_d_out_27_b),
    .io_d_out_27_valid_b(array_5_io_d_out_27_valid_b),
    .io_d_out_28_a(array_5_io_d_out_28_a),
    .io_d_out_28_valid_a(array_5_io_d_out_28_valid_a),
    .io_d_out_28_b(array_5_io_d_out_28_b),
    .io_d_out_28_valid_b(array_5_io_d_out_28_valid_b),
    .io_d_out_29_a(array_5_io_d_out_29_a),
    .io_d_out_29_valid_a(array_5_io_d_out_29_valid_a),
    .io_d_out_29_b(array_5_io_d_out_29_b),
    .io_d_out_29_valid_b(array_5_io_d_out_29_valid_b),
    .io_d_out_30_a(array_5_io_d_out_30_a),
    .io_d_out_30_valid_a(array_5_io_d_out_30_valid_a),
    .io_d_out_30_b(array_5_io_d_out_30_b),
    .io_d_out_30_valid_b(array_5_io_d_out_30_valid_b),
    .io_d_out_31_a(array_5_io_d_out_31_a),
    .io_d_out_31_valid_a(array_5_io_d_out_31_valid_a),
    .io_d_out_31_b(array_5_io_d_out_31_b),
    .io_d_out_31_valid_b(array_5_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_5_io_wr_en_mem1),
    .io_wr_en_mem2(array_5_io_wr_en_mem2),
    .io_wr_en_mem3(array_5_io_wr_en_mem3),
    .io_wr_en_mem4(array_5_io_wr_en_mem4),
    .io_wr_en_mem5(array_5_io_wr_en_mem5),
    .io_wr_en_mem6(array_5_io_wr_en_mem6),
    .io_wr_instr_mem1(array_5_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_5_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_5_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_5_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_5_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_5_io_wr_instr_mem6),
    .io_PC1_in(array_5_io_PC1_in),
    .io_PC6_out(array_5_io_PC6_out),
    .io_Addr_in(array_5_io_Addr_in),
    .io_Addr_out(array_5_io_Addr_out),
    .io_Tag_in_Tag(array_5_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_5_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_5_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_5_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_6 ( // @[Array.scala 41:54]
    .clock(array_6_clock),
    .reset(array_6_reset),
    .io_d_in_0_a(array_6_io_d_in_0_a),
    .io_d_in_0_valid_a(array_6_io_d_in_0_valid_a),
    .io_d_in_0_b(array_6_io_d_in_0_b),
    .io_d_in_1_a(array_6_io_d_in_1_a),
    .io_d_in_1_valid_a(array_6_io_d_in_1_valid_a),
    .io_d_in_1_b(array_6_io_d_in_1_b),
    .io_d_in_2_a(array_6_io_d_in_2_a),
    .io_d_in_2_valid_a(array_6_io_d_in_2_valid_a),
    .io_d_in_2_b(array_6_io_d_in_2_b),
    .io_d_in_3_a(array_6_io_d_in_3_a),
    .io_d_in_3_valid_a(array_6_io_d_in_3_valid_a),
    .io_d_in_3_b(array_6_io_d_in_3_b),
    .io_d_in_4_a(array_6_io_d_in_4_a),
    .io_d_in_4_valid_a(array_6_io_d_in_4_valid_a),
    .io_d_in_4_b(array_6_io_d_in_4_b),
    .io_d_in_5_a(array_6_io_d_in_5_a),
    .io_d_in_5_valid_a(array_6_io_d_in_5_valid_a),
    .io_d_in_5_b(array_6_io_d_in_5_b),
    .io_d_in_6_a(array_6_io_d_in_6_a),
    .io_d_in_6_valid_a(array_6_io_d_in_6_valid_a),
    .io_d_in_6_b(array_6_io_d_in_6_b),
    .io_d_in_7_a(array_6_io_d_in_7_a),
    .io_d_in_7_valid_a(array_6_io_d_in_7_valid_a),
    .io_d_in_7_b(array_6_io_d_in_7_b),
    .io_d_in_8_a(array_6_io_d_in_8_a),
    .io_d_in_8_valid_a(array_6_io_d_in_8_valid_a),
    .io_d_in_8_b(array_6_io_d_in_8_b),
    .io_d_in_9_a(array_6_io_d_in_9_a),
    .io_d_in_9_valid_a(array_6_io_d_in_9_valid_a),
    .io_d_in_9_b(array_6_io_d_in_9_b),
    .io_d_in_10_a(array_6_io_d_in_10_a),
    .io_d_in_10_valid_a(array_6_io_d_in_10_valid_a),
    .io_d_in_10_b(array_6_io_d_in_10_b),
    .io_d_in_11_a(array_6_io_d_in_11_a),
    .io_d_in_11_valid_a(array_6_io_d_in_11_valid_a),
    .io_d_in_11_b(array_6_io_d_in_11_b),
    .io_d_in_12_a(array_6_io_d_in_12_a),
    .io_d_in_12_valid_a(array_6_io_d_in_12_valid_a),
    .io_d_in_12_b(array_6_io_d_in_12_b),
    .io_d_in_13_a(array_6_io_d_in_13_a),
    .io_d_in_13_valid_a(array_6_io_d_in_13_valid_a),
    .io_d_in_13_b(array_6_io_d_in_13_b),
    .io_d_in_14_a(array_6_io_d_in_14_a),
    .io_d_in_14_valid_a(array_6_io_d_in_14_valid_a),
    .io_d_in_14_b(array_6_io_d_in_14_b),
    .io_d_in_15_a(array_6_io_d_in_15_a),
    .io_d_in_15_valid_a(array_6_io_d_in_15_valid_a),
    .io_d_in_15_b(array_6_io_d_in_15_b),
    .io_d_in_16_a(array_6_io_d_in_16_a),
    .io_d_in_16_valid_a(array_6_io_d_in_16_valid_a),
    .io_d_in_16_b(array_6_io_d_in_16_b),
    .io_d_in_17_a(array_6_io_d_in_17_a),
    .io_d_in_17_valid_a(array_6_io_d_in_17_valid_a),
    .io_d_in_17_b(array_6_io_d_in_17_b),
    .io_d_in_18_a(array_6_io_d_in_18_a),
    .io_d_in_18_valid_a(array_6_io_d_in_18_valid_a),
    .io_d_in_18_b(array_6_io_d_in_18_b),
    .io_d_in_19_a(array_6_io_d_in_19_a),
    .io_d_in_19_valid_a(array_6_io_d_in_19_valid_a),
    .io_d_in_19_b(array_6_io_d_in_19_b),
    .io_d_in_20_a(array_6_io_d_in_20_a),
    .io_d_in_20_valid_a(array_6_io_d_in_20_valid_a),
    .io_d_in_20_b(array_6_io_d_in_20_b),
    .io_d_in_21_a(array_6_io_d_in_21_a),
    .io_d_in_21_valid_a(array_6_io_d_in_21_valid_a),
    .io_d_in_21_b(array_6_io_d_in_21_b),
    .io_d_in_22_a(array_6_io_d_in_22_a),
    .io_d_in_22_valid_a(array_6_io_d_in_22_valid_a),
    .io_d_in_22_b(array_6_io_d_in_22_b),
    .io_d_in_23_a(array_6_io_d_in_23_a),
    .io_d_in_23_valid_a(array_6_io_d_in_23_valid_a),
    .io_d_in_23_b(array_6_io_d_in_23_b),
    .io_d_in_24_a(array_6_io_d_in_24_a),
    .io_d_in_24_valid_a(array_6_io_d_in_24_valid_a),
    .io_d_in_24_b(array_6_io_d_in_24_b),
    .io_d_in_25_a(array_6_io_d_in_25_a),
    .io_d_in_25_valid_a(array_6_io_d_in_25_valid_a),
    .io_d_in_25_b(array_6_io_d_in_25_b),
    .io_d_in_26_a(array_6_io_d_in_26_a),
    .io_d_in_26_valid_a(array_6_io_d_in_26_valid_a),
    .io_d_in_26_b(array_6_io_d_in_26_b),
    .io_d_in_27_a(array_6_io_d_in_27_a),
    .io_d_in_27_valid_a(array_6_io_d_in_27_valid_a),
    .io_d_in_27_b(array_6_io_d_in_27_b),
    .io_d_in_28_a(array_6_io_d_in_28_a),
    .io_d_in_28_valid_a(array_6_io_d_in_28_valid_a),
    .io_d_in_28_b(array_6_io_d_in_28_b),
    .io_d_in_29_a(array_6_io_d_in_29_a),
    .io_d_in_29_valid_a(array_6_io_d_in_29_valid_a),
    .io_d_in_29_b(array_6_io_d_in_29_b),
    .io_d_in_30_a(array_6_io_d_in_30_a),
    .io_d_in_30_valid_a(array_6_io_d_in_30_valid_a),
    .io_d_in_30_b(array_6_io_d_in_30_b),
    .io_d_in_31_a(array_6_io_d_in_31_a),
    .io_d_in_31_valid_a(array_6_io_d_in_31_valid_a),
    .io_d_in_31_b(array_6_io_d_in_31_b),
    .io_d_out_0_a(array_6_io_d_out_0_a),
    .io_d_out_0_valid_a(array_6_io_d_out_0_valid_a),
    .io_d_out_0_b(array_6_io_d_out_0_b),
    .io_d_out_0_valid_b(array_6_io_d_out_0_valid_b),
    .io_d_out_1_a(array_6_io_d_out_1_a),
    .io_d_out_1_valid_a(array_6_io_d_out_1_valid_a),
    .io_d_out_1_b(array_6_io_d_out_1_b),
    .io_d_out_1_valid_b(array_6_io_d_out_1_valid_b),
    .io_d_out_2_a(array_6_io_d_out_2_a),
    .io_d_out_2_valid_a(array_6_io_d_out_2_valid_a),
    .io_d_out_2_b(array_6_io_d_out_2_b),
    .io_d_out_2_valid_b(array_6_io_d_out_2_valid_b),
    .io_d_out_3_a(array_6_io_d_out_3_a),
    .io_d_out_3_valid_a(array_6_io_d_out_3_valid_a),
    .io_d_out_3_b(array_6_io_d_out_3_b),
    .io_d_out_3_valid_b(array_6_io_d_out_3_valid_b),
    .io_d_out_4_a(array_6_io_d_out_4_a),
    .io_d_out_4_valid_a(array_6_io_d_out_4_valid_a),
    .io_d_out_4_b(array_6_io_d_out_4_b),
    .io_d_out_4_valid_b(array_6_io_d_out_4_valid_b),
    .io_d_out_5_a(array_6_io_d_out_5_a),
    .io_d_out_5_valid_a(array_6_io_d_out_5_valid_a),
    .io_d_out_5_b(array_6_io_d_out_5_b),
    .io_d_out_5_valid_b(array_6_io_d_out_5_valid_b),
    .io_d_out_6_a(array_6_io_d_out_6_a),
    .io_d_out_6_valid_a(array_6_io_d_out_6_valid_a),
    .io_d_out_6_b(array_6_io_d_out_6_b),
    .io_d_out_6_valid_b(array_6_io_d_out_6_valid_b),
    .io_d_out_7_a(array_6_io_d_out_7_a),
    .io_d_out_7_valid_a(array_6_io_d_out_7_valid_a),
    .io_d_out_7_b(array_6_io_d_out_7_b),
    .io_d_out_7_valid_b(array_6_io_d_out_7_valid_b),
    .io_d_out_8_a(array_6_io_d_out_8_a),
    .io_d_out_8_valid_a(array_6_io_d_out_8_valid_a),
    .io_d_out_8_b(array_6_io_d_out_8_b),
    .io_d_out_8_valid_b(array_6_io_d_out_8_valid_b),
    .io_d_out_9_a(array_6_io_d_out_9_a),
    .io_d_out_9_valid_a(array_6_io_d_out_9_valid_a),
    .io_d_out_9_b(array_6_io_d_out_9_b),
    .io_d_out_9_valid_b(array_6_io_d_out_9_valid_b),
    .io_d_out_10_a(array_6_io_d_out_10_a),
    .io_d_out_10_valid_a(array_6_io_d_out_10_valid_a),
    .io_d_out_10_b(array_6_io_d_out_10_b),
    .io_d_out_10_valid_b(array_6_io_d_out_10_valid_b),
    .io_d_out_11_a(array_6_io_d_out_11_a),
    .io_d_out_11_valid_a(array_6_io_d_out_11_valid_a),
    .io_d_out_11_b(array_6_io_d_out_11_b),
    .io_d_out_11_valid_b(array_6_io_d_out_11_valid_b),
    .io_d_out_12_a(array_6_io_d_out_12_a),
    .io_d_out_12_valid_a(array_6_io_d_out_12_valid_a),
    .io_d_out_12_b(array_6_io_d_out_12_b),
    .io_d_out_12_valid_b(array_6_io_d_out_12_valid_b),
    .io_d_out_13_a(array_6_io_d_out_13_a),
    .io_d_out_13_valid_a(array_6_io_d_out_13_valid_a),
    .io_d_out_13_b(array_6_io_d_out_13_b),
    .io_d_out_13_valid_b(array_6_io_d_out_13_valid_b),
    .io_d_out_14_a(array_6_io_d_out_14_a),
    .io_d_out_14_valid_a(array_6_io_d_out_14_valid_a),
    .io_d_out_14_b(array_6_io_d_out_14_b),
    .io_d_out_14_valid_b(array_6_io_d_out_14_valid_b),
    .io_d_out_15_a(array_6_io_d_out_15_a),
    .io_d_out_15_valid_a(array_6_io_d_out_15_valid_a),
    .io_d_out_15_b(array_6_io_d_out_15_b),
    .io_d_out_15_valid_b(array_6_io_d_out_15_valid_b),
    .io_d_out_16_a(array_6_io_d_out_16_a),
    .io_d_out_16_valid_a(array_6_io_d_out_16_valid_a),
    .io_d_out_16_b(array_6_io_d_out_16_b),
    .io_d_out_16_valid_b(array_6_io_d_out_16_valid_b),
    .io_d_out_17_a(array_6_io_d_out_17_a),
    .io_d_out_17_valid_a(array_6_io_d_out_17_valid_a),
    .io_d_out_17_b(array_6_io_d_out_17_b),
    .io_d_out_17_valid_b(array_6_io_d_out_17_valid_b),
    .io_d_out_18_a(array_6_io_d_out_18_a),
    .io_d_out_18_valid_a(array_6_io_d_out_18_valid_a),
    .io_d_out_18_b(array_6_io_d_out_18_b),
    .io_d_out_18_valid_b(array_6_io_d_out_18_valid_b),
    .io_d_out_19_a(array_6_io_d_out_19_a),
    .io_d_out_19_valid_a(array_6_io_d_out_19_valid_a),
    .io_d_out_19_b(array_6_io_d_out_19_b),
    .io_d_out_19_valid_b(array_6_io_d_out_19_valid_b),
    .io_d_out_20_a(array_6_io_d_out_20_a),
    .io_d_out_20_valid_a(array_6_io_d_out_20_valid_a),
    .io_d_out_20_b(array_6_io_d_out_20_b),
    .io_d_out_20_valid_b(array_6_io_d_out_20_valid_b),
    .io_d_out_21_a(array_6_io_d_out_21_a),
    .io_d_out_21_valid_a(array_6_io_d_out_21_valid_a),
    .io_d_out_21_b(array_6_io_d_out_21_b),
    .io_d_out_21_valid_b(array_6_io_d_out_21_valid_b),
    .io_d_out_22_a(array_6_io_d_out_22_a),
    .io_d_out_22_valid_a(array_6_io_d_out_22_valid_a),
    .io_d_out_22_b(array_6_io_d_out_22_b),
    .io_d_out_22_valid_b(array_6_io_d_out_22_valid_b),
    .io_d_out_23_a(array_6_io_d_out_23_a),
    .io_d_out_23_valid_a(array_6_io_d_out_23_valid_a),
    .io_d_out_23_b(array_6_io_d_out_23_b),
    .io_d_out_23_valid_b(array_6_io_d_out_23_valid_b),
    .io_d_out_24_a(array_6_io_d_out_24_a),
    .io_d_out_24_valid_a(array_6_io_d_out_24_valid_a),
    .io_d_out_24_b(array_6_io_d_out_24_b),
    .io_d_out_24_valid_b(array_6_io_d_out_24_valid_b),
    .io_d_out_25_a(array_6_io_d_out_25_a),
    .io_d_out_25_valid_a(array_6_io_d_out_25_valid_a),
    .io_d_out_25_b(array_6_io_d_out_25_b),
    .io_d_out_25_valid_b(array_6_io_d_out_25_valid_b),
    .io_d_out_26_a(array_6_io_d_out_26_a),
    .io_d_out_26_valid_a(array_6_io_d_out_26_valid_a),
    .io_d_out_26_b(array_6_io_d_out_26_b),
    .io_d_out_26_valid_b(array_6_io_d_out_26_valid_b),
    .io_d_out_27_a(array_6_io_d_out_27_a),
    .io_d_out_27_valid_a(array_6_io_d_out_27_valid_a),
    .io_d_out_27_b(array_6_io_d_out_27_b),
    .io_d_out_27_valid_b(array_6_io_d_out_27_valid_b),
    .io_d_out_28_a(array_6_io_d_out_28_a),
    .io_d_out_28_valid_a(array_6_io_d_out_28_valid_a),
    .io_d_out_28_b(array_6_io_d_out_28_b),
    .io_d_out_28_valid_b(array_6_io_d_out_28_valid_b),
    .io_d_out_29_a(array_6_io_d_out_29_a),
    .io_d_out_29_valid_a(array_6_io_d_out_29_valid_a),
    .io_d_out_29_b(array_6_io_d_out_29_b),
    .io_d_out_29_valid_b(array_6_io_d_out_29_valid_b),
    .io_d_out_30_a(array_6_io_d_out_30_a),
    .io_d_out_30_valid_a(array_6_io_d_out_30_valid_a),
    .io_d_out_30_b(array_6_io_d_out_30_b),
    .io_d_out_30_valid_b(array_6_io_d_out_30_valid_b),
    .io_d_out_31_a(array_6_io_d_out_31_a),
    .io_d_out_31_valid_a(array_6_io_d_out_31_valid_a),
    .io_d_out_31_b(array_6_io_d_out_31_b),
    .io_d_out_31_valid_b(array_6_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_6_io_wr_en_mem1),
    .io_wr_en_mem2(array_6_io_wr_en_mem2),
    .io_wr_en_mem3(array_6_io_wr_en_mem3),
    .io_wr_en_mem4(array_6_io_wr_en_mem4),
    .io_wr_en_mem5(array_6_io_wr_en_mem5),
    .io_wr_en_mem6(array_6_io_wr_en_mem6),
    .io_wr_instr_mem1(array_6_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_6_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_6_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_6_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_6_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_6_io_wr_instr_mem6),
    .io_PC1_in(array_6_io_PC1_in),
    .io_PC6_out(array_6_io_PC6_out),
    .io_Addr_in(array_6_io_Addr_in),
    .io_Addr_out(array_6_io_Addr_out),
    .io_Tag_in_Tag(array_6_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_6_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_6_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_6_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_7 ( // @[Array.scala 41:54]
    .clock(array_7_clock),
    .reset(array_7_reset),
    .io_d_in_0_a(array_7_io_d_in_0_a),
    .io_d_in_0_valid_a(array_7_io_d_in_0_valid_a),
    .io_d_in_0_b(array_7_io_d_in_0_b),
    .io_d_in_1_a(array_7_io_d_in_1_a),
    .io_d_in_1_valid_a(array_7_io_d_in_1_valid_a),
    .io_d_in_1_b(array_7_io_d_in_1_b),
    .io_d_in_2_a(array_7_io_d_in_2_a),
    .io_d_in_2_valid_a(array_7_io_d_in_2_valid_a),
    .io_d_in_2_b(array_7_io_d_in_2_b),
    .io_d_in_3_a(array_7_io_d_in_3_a),
    .io_d_in_3_valid_a(array_7_io_d_in_3_valid_a),
    .io_d_in_3_b(array_7_io_d_in_3_b),
    .io_d_in_4_a(array_7_io_d_in_4_a),
    .io_d_in_4_valid_a(array_7_io_d_in_4_valid_a),
    .io_d_in_4_b(array_7_io_d_in_4_b),
    .io_d_in_5_a(array_7_io_d_in_5_a),
    .io_d_in_5_valid_a(array_7_io_d_in_5_valid_a),
    .io_d_in_5_b(array_7_io_d_in_5_b),
    .io_d_in_6_a(array_7_io_d_in_6_a),
    .io_d_in_6_valid_a(array_7_io_d_in_6_valid_a),
    .io_d_in_6_b(array_7_io_d_in_6_b),
    .io_d_in_7_a(array_7_io_d_in_7_a),
    .io_d_in_7_valid_a(array_7_io_d_in_7_valid_a),
    .io_d_in_7_b(array_7_io_d_in_7_b),
    .io_d_in_8_a(array_7_io_d_in_8_a),
    .io_d_in_8_valid_a(array_7_io_d_in_8_valid_a),
    .io_d_in_8_b(array_7_io_d_in_8_b),
    .io_d_in_9_a(array_7_io_d_in_9_a),
    .io_d_in_9_valid_a(array_7_io_d_in_9_valid_a),
    .io_d_in_9_b(array_7_io_d_in_9_b),
    .io_d_in_10_a(array_7_io_d_in_10_a),
    .io_d_in_10_valid_a(array_7_io_d_in_10_valid_a),
    .io_d_in_10_b(array_7_io_d_in_10_b),
    .io_d_in_11_a(array_7_io_d_in_11_a),
    .io_d_in_11_valid_a(array_7_io_d_in_11_valid_a),
    .io_d_in_11_b(array_7_io_d_in_11_b),
    .io_d_in_12_a(array_7_io_d_in_12_a),
    .io_d_in_12_valid_a(array_7_io_d_in_12_valid_a),
    .io_d_in_12_b(array_7_io_d_in_12_b),
    .io_d_in_13_a(array_7_io_d_in_13_a),
    .io_d_in_13_valid_a(array_7_io_d_in_13_valid_a),
    .io_d_in_13_b(array_7_io_d_in_13_b),
    .io_d_in_14_a(array_7_io_d_in_14_a),
    .io_d_in_14_valid_a(array_7_io_d_in_14_valid_a),
    .io_d_in_14_b(array_7_io_d_in_14_b),
    .io_d_in_15_a(array_7_io_d_in_15_a),
    .io_d_in_15_valid_a(array_7_io_d_in_15_valid_a),
    .io_d_in_15_b(array_7_io_d_in_15_b),
    .io_d_in_16_a(array_7_io_d_in_16_a),
    .io_d_in_16_valid_a(array_7_io_d_in_16_valid_a),
    .io_d_in_16_b(array_7_io_d_in_16_b),
    .io_d_in_17_a(array_7_io_d_in_17_a),
    .io_d_in_17_valid_a(array_7_io_d_in_17_valid_a),
    .io_d_in_17_b(array_7_io_d_in_17_b),
    .io_d_in_18_a(array_7_io_d_in_18_a),
    .io_d_in_18_valid_a(array_7_io_d_in_18_valid_a),
    .io_d_in_18_b(array_7_io_d_in_18_b),
    .io_d_in_19_a(array_7_io_d_in_19_a),
    .io_d_in_19_valid_a(array_7_io_d_in_19_valid_a),
    .io_d_in_19_b(array_7_io_d_in_19_b),
    .io_d_in_20_a(array_7_io_d_in_20_a),
    .io_d_in_20_valid_a(array_7_io_d_in_20_valid_a),
    .io_d_in_20_b(array_7_io_d_in_20_b),
    .io_d_in_21_a(array_7_io_d_in_21_a),
    .io_d_in_21_valid_a(array_7_io_d_in_21_valid_a),
    .io_d_in_21_b(array_7_io_d_in_21_b),
    .io_d_in_22_a(array_7_io_d_in_22_a),
    .io_d_in_22_valid_a(array_7_io_d_in_22_valid_a),
    .io_d_in_22_b(array_7_io_d_in_22_b),
    .io_d_in_23_a(array_7_io_d_in_23_a),
    .io_d_in_23_valid_a(array_7_io_d_in_23_valid_a),
    .io_d_in_23_b(array_7_io_d_in_23_b),
    .io_d_in_24_a(array_7_io_d_in_24_a),
    .io_d_in_24_valid_a(array_7_io_d_in_24_valid_a),
    .io_d_in_24_b(array_7_io_d_in_24_b),
    .io_d_in_25_a(array_7_io_d_in_25_a),
    .io_d_in_25_valid_a(array_7_io_d_in_25_valid_a),
    .io_d_in_25_b(array_7_io_d_in_25_b),
    .io_d_in_26_a(array_7_io_d_in_26_a),
    .io_d_in_26_valid_a(array_7_io_d_in_26_valid_a),
    .io_d_in_26_b(array_7_io_d_in_26_b),
    .io_d_in_27_a(array_7_io_d_in_27_a),
    .io_d_in_27_valid_a(array_7_io_d_in_27_valid_a),
    .io_d_in_27_b(array_7_io_d_in_27_b),
    .io_d_in_28_a(array_7_io_d_in_28_a),
    .io_d_in_28_valid_a(array_7_io_d_in_28_valid_a),
    .io_d_in_28_b(array_7_io_d_in_28_b),
    .io_d_in_29_a(array_7_io_d_in_29_a),
    .io_d_in_29_valid_a(array_7_io_d_in_29_valid_a),
    .io_d_in_29_b(array_7_io_d_in_29_b),
    .io_d_in_30_a(array_7_io_d_in_30_a),
    .io_d_in_30_valid_a(array_7_io_d_in_30_valid_a),
    .io_d_in_30_b(array_7_io_d_in_30_b),
    .io_d_in_31_a(array_7_io_d_in_31_a),
    .io_d_in_31_valid_a(array_7_io_d_in_31_valid_a),
    .io_d_in_31_b(array_7_io_d_in_31_b),
    .io_d_out_0_a(array_7_io_d_out_0_a),
    .io_d_out_0_valid_a(array_7_io_d_out_0_valid_a),
    .io_d_out_0_b(array_7_io_d_out_0_b),
    .io_d_out_0_valid_b(array_7_io_d_out_0_valid_b),
    .io_d_out_1_a(array_7_io_d_out_1_a),
    .io_d_out_1_valid_a(array_7_io_d_out_1_valid_a),
    .io_d_out_1_b(array_7_io_d_out_1_b),
    .io_d_out_1_valid_b(array_7_io_d_out_1_valid_b),
    .io_d_out_2_a(array_7_io_d_out_2_a),
    .io_d_out_2_valid_a(array_7_io_d_out_2_valid_a),
    .io_d_out_2_b(array_7_io_d_out_2_b),
    .io_d_out_2_valid_b(array_7_io_d_out_2_valid_b),
    .io_d_out_3_a(array_7_io_d_out_3_a),
    .io_d_out_3_valid_a(array_7_io_d_out_3_valid_a),
    .io_d_out_3_b(array_7_io_d_out_3_b),
    .io_d_out_3_valid_b(array_7_io_d_out_3_valid_b),
    .io_d_out_4_a(array_7_io_d_out_4_a),
    .io_d_out_4_valid_a(array_7_io_d_out_4_valid_a),
    .io_d_out_4_b(array_7_io_d_out_4_b),
    .io_d_out_4_valid_b(array_7_io_d_out_4_valid_b),
    .io_d_out_5_a(array_7_io_d_out_5_a),
    .io_d_out_5_valid_a(array_7_io_d_out_5_valid_a),
    .io_d_out_5_b(array_7_io_d_out_5_b),
    .io_d_out_5_valid_b(array_7_io_d_out_5_valid_b),
    .io_d_out_6_a(array_7_io_d_out_6_a),
    .io_d_out_6_valid_a(array_7_io_d_out_6_valid_a),
    .io_d_out_6_b(array_7_io_d_out_6_b),
    .io_d_out_6_valid_b(array_7_io_d_out_6_valid_b),
    .io_d_out_7_a(array_7_io_d_out_7_a),
    .io_d_out_7_valid_a(array_7_io_d_out_7_valid_a),
    .io_d_out_7_b(array_7_io_d_out_7_b),
    .io_d_out_7_valid_b(array_7_io_d_out_7_valid_b),
    .io_d_out_8_a(array_7_io_d_out_8_a),
    .io_d_out_8_valid_a(array_7_io_d_out_8_valid_a),
    .io_d_out_8_b(array_7_io_d_out_8_b),
    .io_d_out_8_valid_b(array_7_io_d_out_8_valid_b),
    .io_d_out_9_a(array_7_io_d_out_9_a),
    .io_d_out_9_valid_a(array_7_io_d_out_9_valid_a),
    .io_d_out_9_b(array_7_io_d_out_9_b),
    .io_d_out_9_valid_b(array_7_io_d_out_9_valid_b),
    .io_d_out_10_a(array_7_io_d_out_10_a),
    .io_d_out_10_valid_a(array_7_io_d_out_10_valid_a),
    .io_d_out_10_b(array_7_io_d_out_10_b),
    .io_d_out_10_valid_b(array_7_io_d_out_10_valid_b),
    .io_d_out_11_a(array_7_io_d_out_11_a),
    .io_d_out_11_valid_a(array_7_io_d_out_11_valid_a),
    .io_d_out_11_b(array_7_io_d_out_11_b),
    .io_d_out_11_valid_b(array_7_io_d_out_11_valid_b),
    .io_d_out_12_a(array_7_io_d_out_12_a),
    .io_d_out_12_valid_a(array_7_io_d_out_12_valid_a),
    .io_d_out_12_b(array_7_io_d_out_12_b),
    .io_d_out_12_valid_b(array_7_io_d_out_12_valid_b),
    .io_d_out_13_a(array_7_io_d_out_13_a),
    .io_d_out_13_valid_a(array_7_io_d_out_13_valid_a),
    .io_d_out_13_b(array_7_io_d_out_13_b),
    .io_d_out_13_valid_b(array_7_io_d_out_13_valid_b),
    .io_d_out_14_a(array_7_io_d_out_14_a),
    .io_d_out_14_valid_a(array_7_io_d_out_14_valid_a),
    .io_d_out_14_b(array_7_io_d_out_14_b),
    .io_d_out_14_valid_b(array_7_io_d_out_14_valid_b),
    .io_d_out_15_a(array_7_io_d_out_15_a),
    .io_d_out_15_valid_a(array_7_io_d_out_15_valid_a),
    .io_d_out_15_b(array_7_io_d_out_15_b),
    .io_d_out_15_valid_b(array_7_io_d_out_15_valid_b),
    .io_d_out_16_a(array_7_io_d_out_16_a),
    .io_d_out_16_valid_a(array_7_io_d_out_16_valid_a),
    .io_d_out_16_b(array_7_io_d_out_16_b),
    .io_d_out_16_valid_b(array_7_io_d_out_16_valid_b),
    .io_d_out_17_a(array_7_io_d_out_17_a),
    .io_d_out_17_valid_a(array_7_io_d_out_17_valid_a),
    .io_d_out_17_b(array_7_io_d_out_17_b),
    .io_d_out_17_valid_b(array_7_io_d_out_17_valid_b),
    .io_d_out_18_a(array_7_io_d_out_18_a),
    .io_d_out_18_valid_a(array_7_io_d_out_18_valid_a),
    .io_d_out_18_b(array_7_io_d_out_18_b),
    .io_d_out_18_valid_b(array_7_io_d_out_18_valid_b),
    .io_d_out_19_a(array_7_io_d_out_19_a),
    .io_d_out_19_valid_a(array_7_io_d_out_19_valid_a),
    .io_d_out_19_b(array_7_io_d_out_19_b),
    .io_d_out_19_valid_b(array_7_io_d_out_19_valid_b),
    .io_d_out_20_a(array_7_io_d_out_20_a),
    .io_d_out_20_valid_a(array_7_io_d_out_20_valid_a),
    .io_d_out_20_b(array_7_io_d_out_20_b),
    .io_d_out_20_valid_b(array_7_io_d_out_20_valid_b),
    .io_d_out_21_a(array_7_io_d_out_21_a),
    .io_d_out_21_valid_a(array_7_io_d_out_21_valid_a),
    .io_d_out_21_b(array_7_io_d_out_21_b),
    .io_d_out_21_valid_b(array_7_io_d_out_21_valid_b),
    .io_d_out_22_a(array_7_io_d_out_22_a),
    .io_d_out_22_valid_a(array_7_io_d_out_22_valid_a),
    .io_d_out_22_b(array_7_io_d_out_22_b),
    .io_d_out_22_valid_b(array_7_io_d_out_22_valid_b),
    .io_d_out_23_a(array_7_io_d_out_23_a),
    .io_d_out_23_valid_a(array_7_io_d_out_23_valid_a),
    .io_d_out_23_b(array_7_io_d_out_23_b),
    .io_d_out_23_valid_b(array_7_io_d_out_23_valid_b),
    .io_d_out_24_a(array_7_io_d_out_24_a),
    .io_d_out_24_valid_a(array_7_io_d_out_24_valid_a),
    .io_d_out_24_b(array_7_io_d_out_24_b),
    .io_d_out_24_valid_b(array_7_io_d_out_24_valid_b),
    .io_d_out_25_a(array_7_io_d_out_25_a),
    .io_d_out_25_valid_a(array_7_io_d_out_25_valid_a),
    .io_d_out_25_b(array_7_io_d_out_25_b),
    .io_d_out_25_valid_b(array_7_io_d_out_25_valid_b),
    .io_d_out_26_a(array_7_io_d_out_26_a),
    .io_d_out_26_valid_a(array_7_io_d_out_26_valid_a),
    .io_d_out_26_b(array_7_io_d_out_26_b),
    .io_d_out_26_valid_b(array_7_io_d_out_26_valid_b),
    .io_d_out_27_a(array_7_io_d_out_27_a),
    .io_d_out_27_valid_a(array_7_io_d_out_27_valid_a),
    .io_d_out_27_b(array_7_io_d_out_27_b),
    .io_d_out_27_valid_b(array_7_io_d_out_27_valid_b),
    .io_d_out_28_a(array_7_io_d_out_28_a),
    .io_d_out_28_valid_a(array_7_io_d_out_28_valid_a),
    .io_d_out_28_b(array_7_io_d_out_28_b),
    .io_d_out_28_valid_b(array_7_io_d_out_28_valid_b),
    .io_d_out_29_a(array_7_io_d_out_29_a),
    .io_d_out_29_valid_a(array_7_io_d_out_29_valid_a),
    .io_d_out_29_b(array_7_io_d_out_29_b),
    .io_d_out_29_valid_b(array_7_io_d_out_29_valid_b),
    .io_d_out_30_a(array_7_io_d_out_30_a),
    .io_d_out_30_valid_a(array_7_io_d_out_30_valid_a),
    .io_d_out_30_b(array_7_io_d_out_30_b),
    .io_d_out_30_valid_b(array_7_io_d_out_30_valid_b),
    .io_d_out_31_a(array_7_io_d_out_31_a),
    .io_d_out_31_valid_a(array_7_io_d_out_31_valid_a),
    .io_d_out_31_b(array_7_io_d_out_31_b),
    .io_d_out_31_valid_b(array_7_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_7_io_wr_en_mem1),
    .io_wr_en_mem2(array_7_io_wr_en_mem2),
    .io_wr_en_mem3(array_7_io_wr_en_mem3),
    .io_wr_en_mem4(array_7_io_wr_en_mem4),
    .io_wr_en_mem5(array_7_io_wr_en_mem5),
    .io_wr_en_mem6(array_7_io_wr_en_mem6),
    .io_wr_instr_mem1(array_7_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_7_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_7_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_7_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_7_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_7_io_wr_instr_mem6),
    .io_PC1_in(array_7_io_PC1_in),
    .io_PC6_out(array_7_io_PC6_out),
    .io_Addr_in(array_7_io_Addr_in),
    .io_Addr_out(array_7_io_Addr_out),
    .io_Tag_in_Tag(array_7_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_7_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_7_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_7_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_8 ( // @[Array.scala 41:54]
    .clock(array_8_clock),
    .reset(array_8_reset),
    .io_d_in_0_a(array_8_io_d_in_0_a),
    .io_d_in_0_valid_a(array_8_io_d_in_0_valid_a),
    .io_d_in_0_b(array_8_io_d_in_0_b),
    .io_d_in_1_a(array_8_io_d_in_1_a),
    .io_d_in_1_valid_a(array_8_io_d_in_1_valid_a),
    .io_d_in_1_b(array_8_io_d_in_1_b),
    .io_d_in_2_a(array_8_io_d_in_2_a),
    .io_d_in_2_valid_a(array_8_io_d_in_2_valid_a),
    .io_d_in_2_b(array_8_io_d_in_2_b),
    .io_d_in_3_a(array_8_io_d_in_3_a),
    .io_d_in_3_valid_a(array_8_io_d_in_3_valid_a),
    .io_d_in_3_b(array_8_io_d_in_3_b),
    .io_d_in_4_a(array_8_io_d_in_4_a),
    .io_d_in_4_valid_a(array_8_io_d_in_4_valid_a),
    .io_d_in_4_b(array_8_io_d_in_4_b),
    .io_d_in_5_a(array_8_io_d_in_5_a),
    .io_d_in_5_valid_a(array_8_io_d_in_5_valid_a),
    .io_d_in_5_b(array_8_io_d_in_5_b),
    .io_d_in_6_a(array_8_io_d_in_6_a),
    .io_d_in_6_valid_a(array_8_io_d_in_6_valid_a),
    .io_d_in_6_b(array_8_io_d_in_6_b),
    .io_d_in_7_a(array_8_io_d_in_7_a),
    .io_d_in_7_valid_a(array_8_io_d_in_7_valid_a),
    .io_d_in_7_b(array_8_io_d_in_7_b),
    .io_d_in_8_a(array_8_io_d_in_8_a),
    .io_d_in_8_valid_a(array_8_io_d_in_8_valid_a),
    .io_d_in_8_b(array_8_io_d_in_8_b),
    .io_d_in_9_a(array_8_io_d_in_9_a),
    .io_d_in_9_valid_a(array_8_io_d_in_9_valid_a),
    .io_d_in_9_b(array_8_io_d_in_9_b),
    .io_d_in_10_a(array_8_io_d_in_10_a),
    .io_d_in_10_valid_a(array_8_io_d_in_10_valid_a),
    .io_d_in_10_b(array_8_io_d_in_10_b),
    .io_d_in_11_a(array_8_io_d_in_11_a),
    .io_d_in_11_valid_a(array_8_io_d_in_11_valid_a),
    .io_d_in_11_b(array_8_io_d_in_11_b),
    .io_d_in_12_a(array_8_io_d_in_12_a),
    .io_d_in_12_valid_a(array_8_io_d_in_12_valid_a),
    .io_d_in_12_b(array_8_io_d_in_12_b),
    .io_d_in_13_a(array_8_io_d_in_13_a),
    .io_d_in_13_valid_a(array_8_io_d_in_13_valid_a),
    .io_d_in_13_b(array_8_io_d_in_13_b),
    .io_d_in_14_a(array_8_io_d_in_14_a),
    .io_d_in_14_valid_a(array_8_io_d_in_14_valid_a),
    .io_d_in_14_b(array_8_io_d_in_14_b),
    .io_d_in_15_a(array_8_io_d_in_15_a),
    .io_d_in_15_valid_a(array_8_io_d_in_15_valid_a),
    .io_d_in_15_b(array_8_io_d_in_15_b),
    .io_d_in_16_a(array_8_io_d_in_16_a),
    .io_d_in_16_valid_a(array_8_io_d_in_16_valid_a),
    .io_d_in_16_b(array_8_io_d_in_16_b),
    .io_d_in_17_a(array_8_io_d_in_17_a),
    .io_d_in_17_valid_a(array_8_io_d_in_17_valid_a),
    .io_d_in_17_b(array_8_io_d_in_17_b),
    .io_d_in_18_a(array_8_io_d_in_18_a),
    .io_d_in_18_valid_a(array_8_io_d_in_18_valid_a),
    .io_d_in_18_b(array_8_io_d_in_18_b),
    .io_d_in_19_a(array_8_io_d_in_19_a),
    .io_d_in_19_valid_a(array_8_io_d_in_19_valid_a),
    .io_d_in_19_b(array_8_io_d_in_19_b),
    .io_d_in_20_a(array_8_io_d_in_20_a),
    .io_d_in_20_valid_a(array_8_io_d_in_20_valid_a),
    .io_d_in_20_b(array_8_io_d_in_20_b),
    .io_d_in_21_a(array_8_io_d_in_21_a),
    .io_d_in_21_valid_a(array_8_io_d_in_21_valid_a),
    .io_d_in_21_b(array_8_io_d_in_21_b),
    .io_d_in_22_a(array_8_io_d_in_22_a),
    .io_d_in_22_valid_a(array_8_io_d_in_22_valid_a),
    .io_d_in_22_b(array_8_io_d_in_22_b),
    .io_d_in_23_a(array_8_io_d_in_23_a),
    .io_d_in_23_valid_a(array_8_io_d_in_23_valid_a),
    .io_d_in_23_b(array_8_io_d_in_23_b),
    .io_d_in_24_a(array_8_io_d_in_24_a),
    .io_d_in_24_valid_a(array_8_io_d_in_24_valid_a),
    .io_d_in_24_b(array_8_io_d_in_24_b),
    .io_d_in_25_a(array_8_io_d_in_25_a),
    .io_d_in_25_valid_a(array_8_io_d_in_25_valid_a),
    .io_d_in_25_b(array_8_io_d_in_25_b),
    .io_d_in_26_a(array_8_io_d_in_26_a),
    .io_d_in_26_valid_a(array_8_io_d_in_26_valid_a),
    .io_d_in_26_b(array_8_io_d_in_26_b),
    .io_d_in_27_a(array_8_io_d_in_27_a),
    .io_d_in_27_valid_a(array_8_io_d_in_27_valid_a),
    .io_d_in_27_b(array_8_io_d_in_27_b),
    .io_d_in_28_a(array_8_io_d_in_28_a),
    .io_d_in_28_valid_a(array_8_io_d_in_28_valid_a),
    .io_d_in_28_b(array_8_io_d_in_28_b),
    .io_d_in_29_a(array_8_io_d_in_29_a),
    .io_d_in_29_valid_a(array_8_io_d_in_29_valid_a),
    .io_d_in_29_b(array_8_io_d_in_29_b),
    .io_d_in_30_a(array_8_io_d_in_30_a),
    .io_d_in_30_valid_a(array_8_io_d_in_30_valid_a),
    .io_d_in_30_b(array_8_io_d_in_30_b),
    .io_d_in_31_a(array_8_io_d_in_31_a),
    .io_d_in_31_valid_a(array_8_io_d_in_31_valid_a),
    .io_d_in_31_b(array_8_io_d_in_31_b),
    .io_d_out_0_a(array_8_io_d_out_0_a),
    .io_d_out_0_valid_a(array_8_io_d_out_0_valid_a),
    .io_d_out_0_b(array_8_io_d_out_0_b),
    .io_d_out_0_valid_b(array_8_io_d_out_0_valid_b),
    .io_d_out_1_a(array_8_io_d_out_1_a),
    .io_d_out_1_valid_a(array_8_io_d_out_1_valid_a),
    .io_d_out_1_b(array_8_io_d_out_1_b),
    .io_d_out_1_valid_b(array_8_io_d_out_1_valid_b),
    .io_d_out_2_a(array_8_io_d_out_2_a),
    .io_d_out_2_valid_a(array_8_io_d_out_2_valid_a),
    .io_d_out_2_b(array_8_io_d_out_2_b),
    .io_d_out_2_valid_b(array_8_io_d_out_2_valid_b),
    .io_d_out_3_a(array_8_io_d_out_3_a),
    .io_d_out_3_valid_a(array_8_io_d_out_3_valid_a),
    .io_d_out_3_b(array_8_io_d_out_3_b),
    .io_d_out_3_valid_b(array_8_io_d_out_3_valid_b),
    .io_d_out_4_a(array_8_io_d_out_4_a),
    .io_d_out_4_valid_a(array_8_io_d_out_4_valid_a),
    .io_d_out_4_b(array_8_io_d_out_4_b),
    .io_d_out_4_valid_b(array_8_io_d_out_4_valid_b),
    .io_d_out_5_a(array_8_io_d_out_5_a),
    .io_d_out_5_valid_a(array_8_io_d_out_5_valid_a),
    .io_d_out_5_b(array_8_io_d_out_5_b),
    .io_d_out_5_valid_b(array_8_io_d_out_5_valid_b),
    .io_d_out_6_a(array_8_io_d_out_6_a),
    .io_d_out_6_valid_a(array_8_io_d_out_6_valid_a),
    .io_d_out_6_b(array_8_io_d_out_6_b),
    .io_d_out_6_valid_b(array_8_io_d_out_6_valid_b),
    .io_d_out_7_a(array_8_io_d_out_7_a),
    .io_d_out_7_valid_a(array_8_io_d_out_7_valid_a),
    .io_d_out_7_b(array_8_io_d_out_7_b),
    .io_d_out_7_valid_b(array_8_io_d_out_7_valid_b),
    .io_d_out_8_a(array_8_io_d_out_8_a),
    .io_d_out_8_valid_a(array_8_io_d_out_8_valid_a),
    .io_d_out_8_b(array_8_io_d_out_8_b),
    .io_d_out_8_valid_b(array_8_io_d_out_8_valid_b),
    .io_d_out_9_a(array_8_io_d_out_9_a),
    .io_d_out_9_valid_a(array_8_io_d_out_9_valid_a),
    .io_d_out_9_b(array_8_io_d_out_9_b),
    .io_d_out_9_valid_b(array_8_io_d_out_9_valid_b),
    .io_d_out_10_a(array_8_io_d_out_10_a),
    .io_d_out_10_valid_a(array_8_io_d_out_10_valid_a),
    .io_d_out_10_b(array_8_io_d_out_10_b),
    .io_d_out_10_valid_b(array_8_io_d_out_10_valid_b),
    .io_d_out_11_a(array_8_io_d_out_11_a),
    .io_d_out_11_valid_a(array_8_io_d_out_11_valid_a),
    .io_d_out_11_b(array_8_io_d_out_11_b),
    .io_d_out_11_valid_b(array_8_io_d_out_11_valid_b),
    .io_d_out_12_a(array_8_io_d_out_12_a),
    .io_d_out_12_valid_a(array_8_io_d_out_12_valid_a),
    .io_d_out_12_b(array_8_io_d_out_12_b),
    .io_d_out_12_valid_b(array_8_io_d_out_12_valid_b),
    .io_d_out_13_a(array_8_io_d_out_13_a),
    .io_d_out_13_valid_a(array_8_io_d_out_13_valid_a),
    .io_d_out_13_b(array_8_io_d_out_13_b),
    .io_d_out_13_valid_b(array_8_io_d_out_13_valid_b),
    .io_d_out_14_a(array_8_io_d_out_14_a),
    .io_d_out_14_valid_a(array_8_io_d_out_14_valid_a),
    .io_d_out_14_b(array_8_io_d_out_14_b),
    .io_d_out_14_valid_b(array_8_io_d_out_14_valid_b),
    .io_d_out_15_a(array_8_io_d_out_15_a),
    .io_d_out_15_valid_a(array_8_io_d_out_15_valid_a),
    .io_d_out_15_b(array_8_io_d_out_15_b),
    .io_d_out_15_valid_b(array_8_io_d_out_15_valid_b),
    .io_d_out_16_a(array_8_io_d_out_16_a),
    .io_d_out_16_valid_a(array_8_io_d_out_16_valid_a),
    .io_d_out_16_b(array_8_io_d_out_16_b),
    .io_d_out_16_valid_b(array_8_io_d_out_16_valid_b),
    .io_d_out_17_a(array_8_io_d_out_17_a),
    .io_d_out_17_valid_a(array_8_io_d_out_17_valid_a),
    .io_d_out_17_b(array_8_io_d_out_17_b),
    .io_d_out_17_valid_b(array_8_io_d_out_17_valid_b),
    .io_d_out_18_a(array_8_io_d_out_18_a),
    .io_d_out_18_valid_a(array_8_io_d_out_18_valid_a),
    .io_d_out_18_b(array_8_io_d_out_18_b),
    .io_d_out_18_valid_b(array_8_io_d_out_18_valid_b),
    .io_d_out_19_a(array_8_io_d_out_19_a),
    .io_d_out_19_valid_a(array_8_io_d_out_19_valid_a),
    .io_d_out_19_b(array_8_io_d_out_19_b),
    .io_d_out_19_valid_b(array_8_io_d_out_19_valid_b),
    .io_d_out_20_a(array_8_io_d_out_20_a),
    .io_d_out_20_valid_a(array_8_io_d_out_20_valid_a),
    .io_d_out_20_b(array_8_io_d_out_20_b),
    .io_d_out_20_valid_b(array_8_io_d_out_20_valid_b),
    .io_d_out_21_a(array_8_io_d_out_21_a),
    .io_d_out_21_valid_a(array_8_io_d_out_21_valid_a),
    .io_d_out_21_b(array_8_io_d_out_21_b),
    .io_d_out_21_valid_b(array_8_io_d_out_21_valid_b),
    .io_d_out_22_a(array_8_io_d_out_22_a),
    .io_d_out_22_valid_a(array_8_io_d_out_22_valid_a),
    .io_d_out_22_b(array_8_io_d_out_22_b),
    .io_d_out_22_valid_b(array_8_io_d_out_22_valid_b),
    .io_d_out_23_a(array_8_io_d_out_23_a),
    .io_d_out_23_valid_a(array_8_io_d_out_23_valid_a),
    .io_d_out_23_b(array_8_io_d_out_23_b),
    .io_d_out_23_valid_b(array_8_io_d_out_23_valid_b),
    .io_d_out_24_a(array_8_io_d_out_24_a),
    .io_d_out_24_valid_a(array_8_io_d_out_24_valid_a),
    .io_d_out_24_b(array_8_io_d_out_24_b),
    .io_d_out_24_valid_b(array_8_io_d_out_24_valid_b),
    .io_d_out_25_a(array_8_io_d_out_25_a),
    .io_d_out_25_valid_a(array_8_io_d_out_25_valid_a),
    .io_d_out_25_b(array_8_io_d_out_25_b),
    .io_d_out_25_valid_b(array_8_io_d_out_25_valid_b),
    .io_d_out_26_a(array_8_io_d_out_26_a),
    .io_d_out_26_valid_a(array_8_io_d_out_26_valid_a),
    .io_d_out_26_b(array_8_io_d_out_26_b),
    .io_d_out_26_valid_b(array_8_io_d_out_26_valid_b),
    .io_d_out_27_a(array_8_io_d_out_27_a),
    .io_d_out_27_valid_a(array_8_io_d_out_27_valid_a),
    .io_d_out_27_b(array_8_io_d_out_27_b),
    .io_d_out_27_valid_b(array_8_io_d_out_27_valid_b),
    .io_d_out_28_a(array_8_io_d_out_28_a),
    .io_d_out_28_valid_a(array_8_io_d_out_28_valid_a),
    .io_d_out_28_b(array_8_io_d_out_28_b),
    .io_d_out_28_valid_b(array_8_io_d_out_28_valid_b),
    .io_d_out_29_a(array_8_io_d_out_29_a),
    .io_d_out_29_valid_a(array_8_io_d_out_29_valid_a),
    .io_d_out_29_b(array_8_io_d_out_29_b),
    .io_d_out_29_valid_b(array_8_io_d_out_29_valid_b),
    .io_d_out_30_a(array_8_io_d_out_30_a),
    .io_d_out_30_valid_a(array_8_io_d_out_30_valid_a),
    .io_d_out_30_b(array_8_io_d_out_30_b),
    .io_d_out_30_valid_b(array_8_io_d_out_30_valid_b),
    .io_d_out_31_a(array_8_io_d_out_31_a),
    .io_d_out_31_valid_a(array_8_io_d_out_31_valid_a),
    .io_d_out_31_b(array_8_io_d_out_31_b),
    .io_d_out_31_valid_b(array_8_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_8_io_wr_en_mem1),
    .io_wr_en_mem2(array_8_io_wr_en_mem2),
    .io_wr_en_mem3(array_8_io_wr_en_mem3),
    .io_wr_en_mem4(array_8_io_wr_en_mem4),
    .io_wr_en_mem5(array_8_io_wr_en_mem5),
    .io_wr_en_mem6(array_8_io_wr_en_mem6),
    .io_wr_instr_mem1(array_8_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_8_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_8_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_8_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_8_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_8_io_wr_instr_mem6),
    .io_PC1_in(array_8_io_PC1_in),
    .io_PC6_out(array_8_io_PC6_out),
    .io_Addr_in(array_8_io_Addr_in),
    .io_Addr_out(array_8_io_Addr_out),
    .io_Tag_in_Tag(array_8_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_8_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_8_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_8_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_9 ( // @[Array.scala 41:54]
    .clock(array_9_clock),
    .reset(array_9_reset),
    .io_d_in_0_a(array_9_io_d_in_0_a),
    .io_d_in_0_valid_a(array_9_io_d_in_0_valid_a),
    .io_d_in_0_b(array_9_io_d_in_0_b),
    .io_d_in_1_a(array_9_io_d_in_1_a),
    .io_d_in_1_valid_a(array_9_io_d_in_1_valid_a),
    .io_d_in_1_b(array_9_io_d_in_1_b),
    .io_d_in_2_a(array_9_io_d_in_2_a),
    .io_d_in_2_valid_a(array_9_io_d_in_2_valid_a),
    .io_d_in_2_b(array_9_io_d_in_2_b),
    .io_d_in_3_a(array_9_io_d_in_3_a),
    .io_d_in_3_valid_a(array_9_io_d_in_3_valid_a),
    .io_d_in_3_b(array_9_io_d_in_3_b),
    .io_d_in_4_a(array_9_io_d_in_4_a),
    .io_d_in_4_valid_a(array_9_io_d_in_4_valid_a),
    .io_d_in_4_b(array_9_io_d_in_4_b),
    .io_d_in_5_a(array_9_io_d_in_5_a),
    .io_d_in_5_valid_a(array_9_io_d_in_5_valid_a),
    .io_d_in_5_b(array_9_io_d_in_5_b),
    .io_d_in_6_a(array_9_io_d_in_6_a),
    .io_d_in_6_valid_a(array_9_io_d_in_6_valid_a),
    .io_d_in_6_b(array_9_io_d_in_6_b),
    .io_d_in_7_a(array_9_io_d_in_7_a),
    .io_d_in_7_valid_a(array_9_io_d_in_7_valid_a),
    .io_d_in_7_b(array_9_io_d_in_7_b),
    .io_d_in_8_a(array_9_io_d_in_8_a),
    .io_d_in_8_valid_a(array_9_io_d_in_8_valid_a),
    .io_d_in_8_b(array_9_io_d_in_8_b),
    .io_d_in_9_a(array_9_io_d_in_9_a),
    .io_d_in_9_valid_a(array_9_io_d_in_9_valid_a),
    .io_d_in_9_b(array_9_io_d_in_9_b),
    .io_d_in_10_a(array_9_io_d_in_10_a),
    .io_d_in_10_valid_a(array_9_io_d_in_10_valid_a),
    .io_d_in_10_b(array_9_io_d_in_10_b),
    .io_d_in_11_a(array_9_io_d_in_11_a),
    .io_d_in_11_valid_a(array_9_io_d_in_11_valid_a),
    .io_d_in_11_b(array_9_io_d_in_11_b),
    .io_d_in_12_a(array_9_io_d_in_12_a),
    .io_d_in_12_valid_a(array_9_io_d_in_12_valid_a),
    .io_d_in_12_b(array_9_io_d_in_12_b),
    .io_d_in_13_a(array_9_io_d_in_13_a),
    .io_d_in_13_valid_a(array_9_io_d_in_13_valid_a),
    .io_d_in_13_b(array_9_io_d_in_13_b),
    .io_d_in_14_a(array_9_io_d_in_14_a),
    .io_d_in_14_valid_a(array_9_io_d_in_14_valid_a),
    .io_d_in_14_b(array_9_io_d_in_14_b),
    .io_d_in_15_a(array_9_io_d_in_15_a),
    .io_d_in_15_valid_a(array_9_io_d_in_15_valid_a),
    .io_d_in_15_b(array_9_io_d_in_15_b),
    .io_d_in_16_a(array_9_io_d_in_16_a),
    .io_d_in_16_valid_a(array_9_io_d_in_16_valid_a),
    .io_d_in_16_b(array_9_io_d_in_16_b),
    .io_d_in_17_a(array_9_io_d_in_17_a),
    .io_d_in_17_valid_a(array_9_io_d_in_17_valid_a),
    .io_d_in_17_b(array_9_io_d_in_17_b),
    .io_d_in_18_a(array_9_io_d_in_18_a),
    .io_d_in_18_valid_a(array_9_io_d_in_18_valid_a),
    .io_d_in_18_b(array_9_io_d_in_18_b),
    .io_d_in_19_a(array_9_io_d_in_19_a),
    .io_d_in_19_valid_a(array_9_io_d_in_19_valid_a),
    .io_d_in_19_b(array_9_io_d_in_19_b),
    .io_d_in_20_a(array_9_io_d_in_20_a),
    .io_d_in_20_valid_a(array_9_io_d_in_20_valid_a),
    .io_d_in_20_b(array_9_io_d_in_20_b),
    .io_d_in_21_a(array_9_io_d_in_21_a),
    .io_d_in_21_valid_a(array_9_io_d_in_21_valid_a),
    .io_d_in_21_b(array_9_io_d_in_21_b),
    .io_d_in_22_a(array_9_io_d_in_22_a),
    .io_d_in_22_valid_a(array_9_io_d_in_22_valid_a),
    .io_d_in_22_b(array_9_io_d_in_22_b),
    .io_d_in_23_a(array_9_io_d_in_23_a),
    .io_d_in_23_valid_a(array_9_io_d_in_23_valid_a),
    .io_d_in_23_b(array_9_io_d_in_23_b),
    .io_d_in_24_a(array_9_io_d_in_24_a),
    .io_d_in_24_valid_a(array_9_io_d_in_24_valid_a),
    .io_d_in_24_b(array_9_io_d_in_24_b),
    .io_d_in_25_a(array_9_io_d_in_25_a),
    .io_d_in_25_valid_a(array_9_io_d_in_25_valid_a),
    .io_d_in_25_b(array_9_io_d_in_25_b),
    .io_d_in_26_a(array_9_io_d_in_26_a),
    .io_d_in_26_valid_a(array_9_io_d_in_26_valid_a),
    .io_d_in_26_b(array_9_io_d_in_26_b),
    .io_d_in_27_a(array_9_io_d_in_27_a),
    .io_d_in_27_valid_a(array_9_io_d_in_27_valid_a),
    .io_d_in_27_b(array_9_io_d_in_27_b),
    .io_d_in_28_a(array_9_io_d_in_28_a),
    .io_d_in_28_valid_a(array_9_io_d_in_28_valid_a),
    .io_d_in_28_b(array_9_io_d_in_28_b),
    .io_d_in_29_a(array_9_io_d_in_29_a),
    .io_d_in_29_valid_a(array_9_io_d_in_29_valid_a),
    .io_d_in_29_b(array_9_io_d_in_29_b),
    .io_d_in_30_a(array_9_io_d_in_30_a),
    .io_d_in_30_valid_a(array_9_io_d_in_30_valid_a),
    .io_d_in_30_b(array_9_io_d_in_30_b),
    .io_d_in_31_a(array_9_io_d_in_31_a),
    .io_d_in_31_valid_a(array_9_io_d_in_31_valid_a),
    .io_d_in_31_b(array_9_io_d_in_31_b),
    .io_d_out_0_a(array_9_io_d_out_0_a),
    .io_d_out_0_valid_a(array_9_io_d_out_0_valid_a),
    .io_d_out_0_b(array_9_io_d_out_0_b),
    .io_d_out_0_valid_b(array_9_io_d_out_0_valid_b),
    .io_d_out_1_a(array_9_io_d_out_1_a),
    .io_d_out_1_valid_a(array_9_io_d_out_1_valid_a),
    .io_d_out_1_b(array_9_io_d_out_1_b),
    .io_d_out_1_valid_b(array_9_io_d_out_1_valid_b),
    .io_d_out_2_a(array_9_io_d_out_2_a),
    .io_d_out_2_valid_a(array_9_io_d_out_2_valid_a),
    .io_d_out_2_b(array_9_io_d_out_2_b),
    .io_d_out_2_valid_b(array_9_io_d_out_2_valid_b),
    .io_d_out_3_a(array_9_io_d_out_3_a),
    .io_d_out_3_valid_a(array_9_io_d_out_3_valid_a),
    .io_d_out_3_b(array_9_io_d_out_3_b),
    .io_d_out_3_valid_b(array_9_io_d_out_3_valid_b),
    .io_d_out_4_a(array_9_io_d_out_4_a),
    .io_d_out_4_valid_a(array_9_io_d_out_4_valid_a),
    .io_d_out_4_b(array_9_io_d_out_4_b),
    .io_d_out_4_valid_b(array_9_io_d_out_4_valid_b),
    .io_d_out_5_a(array_9_io_d_out_5_a),
    .io_d_out_5_valid_a(array_9_io_d_out_5_valid_a),
    .io_d_out_5_b(array_9_io_d_out_5_b),
    .io_d_out_5_valid_b(array_9_io_d_out_5_valid_b),
    .io_d_out_6_a(array_9_io_d_out_6_a),
    .io_d_out_6_valid_a(array_9_io_d_out_6_valid_a),
    .io_d_out_6_b(array_9_io_d_out_6_b),
    .io_d_out_6_valid_b(array_9_io_d_out_6_valid_b),
    .io_d_out_7_a(array_9_io_d_out_7_a),
    .io_d_out_7_valid_a(array_9_io_d_out_7_valid_a),
    .io_d_out_7_b(array_9_io_d_out_7_b),
    .io_d_out_7_valid_b(array_9_io_d_out_7_valid_b),
    .io_d_out_8_a(array_9_io_d_out_8_a),
    .io_d_out_8_valid_a(array_9_io_d_out_8_valid_a),
    .io_d_out_8_b(array_9_io_d_out_8_b),
    .io_d_out_8_valid_b(array_9_io_d_out_8_valid_b),
    .io_d_out_9_a(array_9_io_d_out_9_a),
    .io_d_out_9_valid_a(array_9_io_d_out_9_valid_a),
    .io_d_out_9_b(array_9_io_d_out_9_b),
    .io_d_out_9_valid_b(array_9_io_d_out_9_valid_b),
    .io_d_out_10_a(array_9_io_d_out_10_a),
    .io_d_out_10_valid_a(array_9_io_d_out_10_valid_a),
    .io_d_out_10_b(array_9_io_d_out_10_b),
    .io_d_out_10_valid_b(array_9_io_d_out_10_valid_b),
    .io_d_out_11_a(array_9_io_d_out_11_a),
    .io_d_out_11_valid_a(array_9_io_d_out_11_valid_a),
    .io_d_out_11_b(array_9_io_d_out_11_b),
    .io_d_out_11_valid_b(array_9_io_d_out_11_valid_b),
    .io_d_out_12_a(array_9_io_d_out_12_a),
    .io_d_out_12_valid_a(array_9_io_d_out_12_valid_a),
    .io_d_out_12_b(array_9_io_d_out_12_b),
    .io_d_out_12_valid_b(array_9_io_d_out_12_valid_b),
    .io_d_out_13_a(array_9_io_d_out_13_a),
    .io_d_out_13_valid_a(array_9_io_d_out_13_valid_a),
    .io_d_out_13_b(array_9_io_d_out_13_b),
    .io_d_out_13_valid_b(array_9_io_d_out_13_valid_b),
    .io_d_out_14_a(array_9_io_d_out_14_a),
    .io_d_out_14_valid_a(array_9_io_d_out_14_valid_a),
    .io_d_out_14_b(array_9_io_d_out_14_b),
    .io_d_out_14_valid_b(array_9_io_d_out_14_valid_b),
    .io_d_out_15_a(array_9_io_d_out_15_a),
    .io_d_out_15_valid_a(array_9_io_d_out_15_valid_a),
    .io_d_out_15_b(array_9_io_d_out_15_b),
    .io_d_out_15_valid_b(array_9_io_d_out_15_valid_b),
    .io_d_out_16_a(array_9_io_d_out_16_a),
    .io_d_out_16_valid_a(array_9_io_d_out_16_valid_a),
    .io_d_out_16_b(array_9_io_d_out_16_b),
    .io_d_out_16_valid_b(array_9_io_d_out_16_valid_b),
    .io_d_out_17_a(array_9_io_d_out_17_a),
    .io_d_out_17_valid_a(array_9_io_d_out_17_valid_a),
    .io_d_out_17_b(array_9_io_d_out_17_b),
    .io_d_out_17_valid_b(array_9_io_d_out_17_valid_b),
    .io_d_out_18_a(array_9_io_d_out_18_a),
    .io_d_out_18_valid_a(array_9_io_d_out_18_valid_a),
    .io_d_out_18_b(array_9_io_d_out_18_b),
    .io_d_out_18_valid_b(array_9_io_d_out_18_valid_b),
    .io_d_out_19_a(array_9_io_d_out_19_a),
    .io_d_out_19_valid_a(array_9_io_d_out_19_valid_a),
    .io_d_out_19_b(array_9_io_d_out_19_b),
    .io_d_out_19_valid_b(array_9_io_d_out_19_valid_b),
    .io_d_out_20_a(array_9_io_d_out_20_a),
    .io_d_out_20_valid_a(array_9_io_d_out_20_valid_a),
    .io_d_out_20_b(array_9_io_d_out_20_b),
    .io_d_out_20_valid_b(array_9_io_d_out_20_valid_b),
    .io_d_out_21_a(array_9_io_d_out_21_a),
    .io_d_out_21_valid_a(array_9_io_d_out_21_valid_a),
    .io_d_out_21_b(array_9_io_d_out_21_b),
    .io_d_out_21_valid_b(array_9_io_d_out_21_valid_b),
    .io_d_out_22_a(array_9_io_d_out_22_a),
    .io_d_out_22_valid_a(array_9_io_d_out_22_valid_a),
    .io_d_out_22_b(array_9_io_d_out_22_b),
    .io_d_out_22_valid_b(array_9_io_d_out_22_valid_b),
    .io_d_out_23_a(array_9_io_d_out_23_a),
    .io_d_out_23_valid_a(array_9_io_d_out_23_valid_a),
    .io_d_out_23_b(array_9_io_d_out_23_b),
    .io_d_out_23_valid_b(array_9_io_d_out_23_valid_b),
    .io_d_out_24_a(array_9_io_d_out_24_a),
    .io_d_out_24_valid_a(array_9_io_d_out_24_valid_a),
    .io_d_out_24_b(array_9_io_d_out_24_b),
    .io_d_out_24_valid_b(array_9_io_d_out_24_valid_b),
    .io_d_out_25_a(array_9_io_d_out_25_a),
    .io_d_out_25_valid_a(array_9_io_d_out_25_valid_a),
    .io_d_out_25_b(array_9_io_d_out_25_b),
    .io_d_out_25_valid_b(array_9_io_d_out_25_valid_b),
    .io_d_out_26_a(array_9_io_d_out_26_a),
    .io_d_out_26_valid_a(array_9_io_d_out_26_valid_a),
    .io_d_out_26_b(array_9_io_d_out_26_b),
    .io_d_out_26_valid_b(array_9_io_d_out_26_valid_b),
    .io_d_out_27_a(array_9_io_d_out_27_a),
    .io_d_out_27_valid_a(array_9_io_d_out_27_valid_a),
    .io_d_out_27_b(array_9_io_d_out_27_b),
    .io_d_out_27_valid_b(array_9_io_d_out_27_valid_b),
    .io_d_out_28_a(array_9_io_d_out_28_a),
    .io_d_out_28_valid_a(array_9_io_d_out_28_valid_a),
    .io_d_out_28_b(array_9_io_d_out_28_b),
    .io_d_out_28_valid_b(array_9_io_d_out_28_valid_b),
    .io_d_out_29_a(array_9_io_d_out_29_a),
    .io_d_out_29_valid_a(array_9_io_d_out_29_valid_a),
    .io_d_out_29_b(array_9_io_d_out_29_b),
    .io_d_out_29_valid_b(array_9_io_d_out_29_valid_b),
    .io_d_out_30_a(array_9_io_d_out_30_a),
    .io_d_out_30_valid_a(array_9_io_d_out_30_valid_a),
    .io_d_out_30_b(array_9_io_d_out_30_b),
    .io_d_out_30_valid_b(array_9_io_d_out_30_valid_b),
    .io_d_out_31_a(array_9_io_d_out_31_a),
    .io_d_out_31_valid_a(array_9_io_d_out_31_valid_a),
    .io_d_out_31_b(array_9_io_d_out_31_b),
    .io_d_out_31_valid_b(array_9_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_9_io_wr_en_mem1),
    .io_wr_en_mem2(array_9_io_wr_en_mem2),
    .io_wr_en_mem3(array_9_io_wr_en_mem3),
    .io_wr_en_mem4(array_9_io_wr_en_mem4),
    .io_wr_en_mem5(array_9_io_wr_en_mem5),
    .io_wr_en_mem6(array_9_io_wr_en_mem6),
    .io_wr_instr_mem1(array_9_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_9_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_9_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_9_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_9_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_9_io_wr_instr_mem6),
    .io_PC1_in(array_9_io_PC1_in),
    .io_PC6_out(array_9_io_PC6_out),
    .io_Addr_in(array_9_io_Addr_in),
    .io_Addr_out(array_9_io_Addr_out),
    .io_Tag_in_Tag(array_9_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_9_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_9_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_9_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_10 ( // @[Array.scala 41:54]
    .clock(array_10_clock),
    .reset(array_10_reset),
    .io_d_in_0_a(array_10_io_d_in_0_a),
    .io_d_in_0_valid_a(array_10_io_d_in_0_valid_a),
    .io_d_in_0_b(array_10_io_d_in_0_b),
    .io_d_in_1_a(array_10_io_d_in_1_a),
    .io_d_in_1_valid_a(array_10_io_d_in_1_valid_a),
    .io_d_in_1_b(array_10_io_d_in_1_b),
    .io_d_in_2_a(array_10_io_d_in_2_a),
    .io_d_in_2_valid_a(array_10_io_d_in_2_valid_a),
    .io_d_in_2_b(array_10_io_d_in_2_b),
    .io_d_in_3_a(array_10_io_d_in_3_a),
    .io_d_in_3_valid_a(array_10_io_d_in_3_valid_a),
    .io_d_in_3_b(array_10_io_d_in_3_b),
    .io_d_in_4_a(array_10_io_d_in_4_a),
    .io_d_in_4_valid_a(array_10_io_d_in_4_valid_a),
    .io_d_in_4_b(array_10_io_d_in_4_b),
    .io_d_in_5_a(array_10_io_d_in_5_a),
    .io_d_in_5_valid_a(array_10_io_d_in_5_valid_a),
    .io_d_in_5_b(array_10_io_d_in_5_b),
    .io_d_in_6_a(array_10_io_d_in_6_a),
    .io_d_in_6_valid_a(array_10_io_d_in_6_valid_a),
    .io_d_in_6_b(array_10_io_d_in_6_b),
    .io_d_in_7_a(array_10_io_d_in_7_a),
    .io_d_in_7_valid_a(array_10_io_d_in_7_valid_a),
    .io_d_in_7_b(array_10_io_d_in_7_b),
    .io_d_in_8_a(array_10_io_d_in_8_a),
    .io_d_in_8_valid_a(array_10_io_d_in_8_valid_a),
    .io_d_in_8_b(array_10_io_d_in_8_b),
    .io_d_in_9_a(array_10_io_d_in_9_a),
    .io_d_in_9_valid_a(array_10_io_d_in_9_valid_a),
    .io_d_in_9_b(array_10_io_d_in_9_b),
    .io_d_in_10_a(array_10_io_d_in_10_a),
    .io_d_in_10_valid_a(array_10_io_d_in_10_valid_a),
    .io_d_in_10_b(array_10_io_d_in_10_b),
    .io_d_in_11_a(array_10_io_d_in_11_a),
    .io_d_in_11_valid_a(array_10_io_d_in_11_valid_a),
    .io_d_in_11_b(array_10_io_d_in_11_b),
    .io_d_in_12_a(array_10_io_d_in_12_a),
    .io_d_in_12_valid_a(array_10_io_d_in_12_valid_a),
    .io_d_in_12_b(array_10_io_d_in_12_b),
    .io_d_in_13_a(array_10_io_d_in_13_a),
    .io_d_in_13_valid_a(array_10_io_d_in_13_valid_a),
    .io_d_in_13_b(array_10_io_d_in_13_b),
    .io_d_in_14_a(array_10_io_d_in_14_a),
    .io_d_in_14_valid_a(array_10_io_d_in_14_valid_a),
    .io_d_in_14_b(array_10_io_d_in_14_b),
    .io_d_in_15_a(array_10_io_d_in_15_a),
    .io_d_in_15_valid_a(array_10_io_d_in_15_valid_a),
    .io_d_in_15_b(array_10_io_d_in_15_b),
    .io_d_in_16_a(array_10_io_d_in_16_a),
    .io_d_in_16_valid_a(array_10_io_d_in_16_valid_a),
    .io_d_in_16_b(array_10_io_d_in_16_b),
    .io_d_in_17_a(array_10_io_d_in_17_a),
    .io_d_in_17_valid_a(array_10_io_d_in_17_valid_a),
    .io_d_in_17_b(array_10_io_d_in_17_b),
    .io_d_in_18_a(array_10_io_d_in_18_a),
    .io_d_in_18_valid_a(array_10_io_d_in_18_valid_a),
    .io_d_in_18_b(array_10_io_d_in_18_b),
    .io_d_in_19_a(array_10_io_d_in_19_a),
    .io_d_in_19_valid_a(array_10_io_d_in_19_valid_a),
    .io_d_in_19_b(array_10_io_d_in_19_b),
    .io_d_in_20_a(array_10_io_d_in_20_a),
    .io_d_in_20_valid_a(array_10_io_d_in_20_valid_a),
    .io_d_in_20_b(array_10_io_d_in_20_b),
    .io_d_in_21_a(array_10_io_d_in_21_a),
    .io_d_in_21_valid_a(array_10_io_d_in_21_valid_a),
    .io_d_in_21_b(array_10_io_d_in_21_b),
    .io_d_in_22_a(array_10_io_d_in_22_a),
    .io_d_in_22_valid_a(array_10_io_d_in_22_valid_a),
    .io_d_in_22_b(array_10_io_d_in_22_b),
    .io_d_in_23_a(array_10_io_d_in_23_a),
    .io_d_in_23_valid_a(array_10_io_d_in_23_valid_a),
    .io_d_in_23_b(array_10_io_d_in_23_b),
    .io_d_in_24_a(array_10_io_d_in_24_a),
    .io_d_in_24_valid_a(array_10_io_d_in_24_valid_a),
    .io_d_in_24_b(array_10_io_d_in_24_b),
    .io_d_in_25_a(array_10_io_d_in_25_a),
    .io_d_in_25_valid_a(array_10_io_d_in_25_valid_a),
    .io_d_in_25_b(array_10_io_d_in_25_b),
    .io_d_in_26_a(array_10_io_d_in_26_a),
    .io_d_in_26_valid_a(array_10_io_d_in_26_valid_a),
    .io_d_in_26_b(array_10_io_d_in_26_b),
    .io_d_in_27_a(array_10_io_d_in_27_a),
    .io_d_in_27_valid_a(array_10_io_d_in_27_valid_a),
    .io_d_in_27_b(array_10_io_d_in_27_b),
    .io_d_in_28_a(array_10_io_d_in_28_a),
    .io_d_in_28_valid_a(array_10_io_d_in_28_valid_a),
    .io_d_in_28_b(array_10_io_d_in_28_b),
    .io_d_in_29_a(array_10_io_d_in_29_a),
    .io_d_in_29_valid_a(array_10_io_d_in_29_valid_a),
    .io_d_in_29_b(array_10_io_d_in_29_b),
    .io_d_in_30_a(array_10_io_d_in_30_a),
    .io_d_in_30_valid_a(array_10_io_d_in_30_valid_a),
    .io_d_in_30_b(array_10_io_d_in_30_b),
    .io_d_in_31_a(array_10_io_d_in_31_a),
    .io_d_in_31_valid_a(array_10_io_d_in_31_valid_a),
    .io_d_in_31_b(array_10_io_d_in_31_b),
    .io_d_out_0_a(array_10_io_d_out_0_a),
    .io_d_out_0_valid_a(array_10_io_d_out_0_valid_a),
    .io_d_out_0_b(array_10_io_d_out_0_b),
    .io_d_out_0_valid_b(array_10_io_d_out_0_valid_b),
    .io_d_out_1_a(array_10_io_d_out_1_a),
    .io_d_out_1_valid_a(array_10_io_d_out_1_valid_a),
    .io_d_out_1_b(array_10_io_d_out_1_b),
    .io_d_out_1_valid_b(array_10_io_d_out_1_valid_b),
    .io_d_out_2_a(array_10_io_d_out_2_a),
    .io_d_out_2_valid_a(array_10_io_d_out_2_valid_a),
    .io_d_out_2_b(array_10_io_d_out_2_b),
    .io_d_out_2_valid_b(array_10_io_d_out_2_valid_b),
    .io_d_out_3_a(array_10_io_d_out_3_a),
    .io_d_out_3_valid_a(array_10_io_d_out_3_valid_a),
    .io_d_out_3_b(array_10_io_d_out_3_b),
    .io_d_out_3_valid_b(array_10_io_d_out_3_valid_b),
    .io_d_out_4_a(array_10_io_d_out_4_a),
    .io_d_out_4_valid_a(array_10_io_d_out_4_valid_a),
    .io_d_out_4_b(array_10_io_d_out_4_b),
    .io_d_out_4_valid_b(array_10_io_d_out_4_valid_b),
    .io_d_out_5_a(array_10_io_d_out_5_a),
    .io_d_out_5_valid_a(array_10_io_d_out_5_valid_a),
    .io_d_out_5_b(array_10_io_d_out_5_b),
    .io_d_out_5_valid_b(array_10_io_d_out_5_valid_b),
    .io_d_out_6_a(array_10_io_d_out_6_a),
    .io_d_out_6_valid_a(array_10_io_d_out_6_valid_a),
    .io_d_out_6_b(array_10_io_d_out_6_b),
    .io_d_out_6_valid_b(array_10_io_d_out_6_valid_b),
    .io_d_out_7_a(array_10_io_d_out_7_a),
    .io_d_out_7_valid_a(array_10_io_d_out_7_valid_a),
    .io_d_out_7_b(array_10_io_d_out_7_b),
    .io_d_out_7_valid_b(array_10_io_d_out_7_valid_b),
    .io_d_out_8_a(array_10_io_d_out_8_a),
    .io_d_out_8_valid_a(array_10_io_d_out_8_valid_a),
    .io_d_out_8_b(array_10_io_d_out_8_b),
    .io_d_out_8_valid_b(array_10_io_d_out_8_valid_b),
    .io_d_out_9_a(array_10_io_d_out_9_a),
    .io_d_out_9_valid_a(array_10_io_d_out_9_valid_a),
    .io_d_out_9_b(array_10_io_d_out_9_b),
    .io_d_out_9_valid_b(array_10_io_d_out_9_valid_b),
    .io_d_out_10_a(array_10_io_d_out_10_a),
    .io_d_out_10_valid_a(array_10_io_d_out_10_valid_a),
    .io_d_out_10_b(array_10_io_d_out_10_b),
    .io_d_out_10_valid_b(array_10_io_d_out_10_valid_b),
    .io_d_out_11_a(array_10_io_d_out_11_a),
    .io_d_out_11_valid_a(array_10_io_d_out_11_valid_a),
    .io_d_out_11_b(array_10_io_d_out_11_b),
    .io_d_out_11_valid_b(array_10_io_d_out_11_valid_b),
    .io_d_out_12_a(array_10_io_d_out_12_a),
    .io_d_out_12_valid_a(array_10_io_d_out_12_valid_a),
    .io_d_out_12_b(array_10_io_d_out_12_b),
    .io_d_out_12_valid_b(array_10_io_d_out_12_valid_b),
    .io_d_out_13_a(array_10_io_d_out_13_a),
    .io_d_out_13_valid_a(array_10_io_d_out_13_valid_a),
    .io_d_out_13_b(array_10_io_d_out_13_b),
    .io_d_out_13_valid_b(array_10_io_d_out_13_valid_b),
    .io_d_out_14_a(array_10_io_d_out_14_a),
    .io_d_out_14_valid_a(array_10_io_d_out_14_valid_a),
    .io_d_out_14_b(array_10_io_d_out_14_b),
    .io_d_out_14_valid_b(array_10_io_d_out_14_valid_b),
    .io_d_out_15_a(array_10_io_d_out_15_a),
    .io_d_out_15_valid_a(array_10_io_d_out_15_valid_a),
    .io_d_out_15_b(array_10_io_d_out_15_b),
    .io_d_out_15_valid_b(array_10_io_d_out_15_valid_b),
    .io_d_out_16_a(array_10_io_d_out_16_a),
    .io_d_out_16_valid_a(array_10_io_d_out_16_valid_a),
    .io_d_out_16_b(array_10_io_d_out_16_b),
    .io_d_out_16_valid_b(array_10_io_d_out_16_valid_b),
    .io_d_out_17_a(array_10_io_d_out_17_a),
    .io_d_out_17_valid_a(array_10_io_d_out_17_valid_a),
    .io_d_out_17_b(array_10_io_d_out_17_b),
    .io_d_out_17_valid_b(array_10_io_d_out_17_valid_b),
    .io_d_out_18_a(array_10_io_d_out_18_a),
    .io_d_out_18_valid_a(array_10_io_d_out_18_valid_a),
    .io_d_out_18_b(array_10_io_d_out_18_b),
    .io_d_out_18_valid_b(array_10_io_d_out_18_valid_b),
    .io_d_out_19_a(array_10_io_d_out_19_a),
    .io_d_out_19_valid_a(array_10_io_d_out_19_valid_a),
    .io_d_out_19_b(array_10_io_d_out_19_b),
    .io_d_out_19_valid_b(array_10_io_d_out_19_valid_b),
    .io_d_out_20_a(array_10_io_d_out_20_a),
    .io_d_out_20_valid_a(array_10_io_d_out_20_valid_a),
    .io_d_out_20_b(array_10_io_d_out_20_b),
    .io_d_out_20_valid_b(array_10_io_d_out_20_valid_b),
    .io_d_out_21_a(array_10_io_d_out_21_a),
    .io_d_out_21_valid_a(array_10_io_d_out_21_valid_a),
    .io_d_out_21_b(array_10_io_d_out_21_b),
    .io_d_out_21_valid_b(array_10_io_d_out_21_valid_b),
    .io_d_out_22_a(array_10_io_d_out_22_a),
    .io_d_out_22_valid_a(array_10_io_d_out_22_valid_a),
    .io_d_out_22_b(array_10_io_d_out_22_b),
    .io_d_out_22_valid_b(array_10_io_d_out_22_valid_b),
    .io_d_out_23_a(array_10_io_d_out_23_a),
    .io_d_out_23_valid_a(array_10_io_d_out_23_valid_a),
    .io_d_out_23_b(array_10_io_d_out_23_b),
    .io_d_out_23_valid_b(array_10_io_d_out_23_valid_b),
    .io_d_out_24_a(array_10_io_d_out_24_a),
    .io_d_out_24_valid_a(array_10_io_d_out_24_valid_a),
    .io_d_out_24_b(array_10_io_d_out_24_b),
    .io_d_out_24_valid_b(array_10_io_d_out_24_valid_b),
    .io_d_out_25_a(array_10_io_d_out_25_a),
    .io_d_out_25_valid_a(array_10_io_d_out_25_valid_a),
    .io_d_out_25_b(array_10_io_d_out_25_b),
    .io_d_out_25_valid_b(array_10_io_d_out_25_valid_b),
    .io_d_out_26_a(array_10_io_d_out_26_a),
    .io_d_out_26_valid_a(array_10_io_d_out_26_valid_a),
    .io_d_out_26_b(array_10_io_d_out_26_b),
    .io_d_out_26_valid_b(array_10_io_d_out_26_valid_b),
    .io_d_out_27_a(array_10_io_d_out_27_a),
    .io_d_out_27_valid_a(array_10_io_d_out_27_valid_a),
    .io_d_out_27_b(array_10_io_d_out_27_b),
    .io_d_out_27_valid_b(array_10_io_d_out_27_valid_b),
    .io_d_out_28_a(array_10_io_d_out_28_a),
    .io_d_out_28_valid_a(array_10_io_d_out_28_valid_a),
    .io_d_out_28_b(array_10_io_d_out_28_b),
    .io_d_out_28_valid_b(array_10_io_d_out_28_valid_b),
    .io_d_out_29_a(array_10_io_d_out_29_a),
    .io_d_out_29_valid_a(array_10_io_d_out_29_valid_a),
    .io_d_out_29_b(array_10_io_d_out_29_b),
    .io_d_out_29_valid_b(array_10_io_d_out_29_valid_b),
    .io_d_out_30_a(array_10_io_d_out_30_a),
    .io_d_out_30_valid_a(array_10_io_d_out_30_valid_a),
    .io_d_out_30_b(array_10_io_d_out_30_b),
    .io_d_out_30_valid_b(array_10_io_d_out_30_valid_b),
    .io_d_out_31_a(array_10_io_d_out_31_a),
    .io_d_out_31_valid_a(array_10_io_d_out_31_valid_a),
    .io_d_out_31_b(array_10_io_d_out_31_b),
    .io_d_out_31_valid_b(array_10_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_10_io_wr_en_mem1),
    .io_wr_en_mem2(array_10_io_wr_en_mem2),
    .io_wr_en_mem3(array_10_io_wr_en_mem3),
    .io_wr_en_mem4(array_10_io_wr_en_mem4),
    .io_wr_en_mem5(array_10_io_wr_en_mem5),
    .io_wr_en_mem6(array_10_io_wr_en_mem6),
    .io_wr_instr_mem1(array_10_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_10_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_10_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_10_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_10_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_10_io_wr_instr_mem6),
    .io_PC1_in(array_10_io_PC1_in),
    .io_PC6_out(array_10_io_PC6_out),
    .io_Addr_in(array_10_io_Addr_in),
    .io_Addr_out(array_10_io_Addr_out),
    .io_Tag_in_Tag(array_10_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_10_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_10_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_10_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_11 ( // @[Array.scala 41:54]
    .clock(array_11_clock),
    .reset(array_11_reset),
    .io_d_in_0_a(array_11_io_d_in_0_a),
    .io_d_in_0_valid_a(array_11_io_d_in_0_valid_a),
    .io_d_in_0_b(array_11_io_d_in_0_b),
    .io_d_in_1_a(array_11_io_d_in_1_a),
    .io_d_in_1_valid_a(array_11_io_d_in_1_valid_a),
    .io_d_in_1_b(array_11_io_d_in_1_b),
    .io_d_in_2_a(array_11_io_d_in_2_a),
    .io_d_in_2_valid_a(array_11_io_d_in_2_valid_a),
    .io_d_in_2_b(array_11_io_d_in_2_b),
    .io_d_in_3_a(array_11_io_d_in_3_a),
    .io_d_in_3_valid_a(array_11_io_d_in_3_valid_a),
    .io_d_in_3_b(array_11_io_d_in_3_b),
    .io_d_in_4_a(array_11_io_d_in_4_a),
    .io_d_in_4_valid_a(array_11_io_d_in_4_valid_a),
    .io_d_in_4_b(array_11_io_d_in_4_b),
    .io_d_in_5_a(array_11_io_d_in_5_a),
    .io_d_in_5_valid_a(array_11_io_d_in_5_valid_a),
    .io_d_in_5_b(array_11_io_d_in_5_b),
    .io_d_in_6_a(array_11_io_d_in_6_a),
    .io_d_in_6_valid_a(array_11_io_d_in_6_valid_a),
    .io_d_in_6_b(array_11_io_d_in_6_b),
    .io_d_in_7_a(array_11_io_d_in_7_a),
    .io_d_in_7_valid_a(array_11_io_d_in_7_valid_a),
    .io_d_in_7_b(array_11_io_d_in_7_b),
    .io_d_in_8_a(array_11_io_d_in_8_a),
    .io_d_in_8_valid_a(array_11_io_d_in_8_valid_a),
    .io_d_in_8_b(array_11_io_d_in_8_b),
    .io_d_in_9_a(array_11_io_d_in_9_a),
    .io_d_in_9_valid_a(array_11_io_d_in_9_valid_a),
    .io_d_in_9_b(array_11_io_d_in_9_b),
    .io_d_in_10_a(array_11_io_d_in_10_a),
    .io_d_in_10_valid_a(array_11_io_d_in_10_valid_a),
    .io_d_in_10_b(array_11_io_d_in_10_b),
    .io_d_in_11_a(array_11_io_d_in_11_a),
    .io_d_in_11_valid_a(array_11_io_d_in_11_valid_a),
    .io_d_in_11_b(array_11_io_d_in_11_b),
    .io_d_in_12_a(array_11_io_d_in_12_a),
    .io_d_in_12_valid_a(array_11_io_d_in_12_valid_a),
    .io_d_in_12_b(array_11_io_d_in_12_b),
    .io_d_in_13_a(array_11_io_d_in_13_a),
    .io_d_in_13_valid_a(array_11_io_d_in_13_valid_a),
    .io_d_in_13_b(array_11_io_d_in_13_b),
    .io_d_in_14_a(array_11_io_d_in_14_a),
    .io_d_in_14_valid_a(array_11_io_d_in_14_valid_a),
    .io_d_in_14_b(array_11_io_d_in_14_b),
    .io_d_in_15_a(array_11_io_d_in_15_a),
    .io_d_in_15_valid_a(array_11_io_d_in_15_valid_a),
    .io_d_in_15_b(array_11_io_d_in_15_b),
    .io_d_in_16_a(array_11_io_d_in_16_a),
    .io_d_in_16_valid_a(array_11_io_d_in_16_valid_a),
    .io_d_in_16_b(array_11_io_d_in_16_b),
    .io_d_in_17_a(array_11_io_d_in_17_a),
    .io_d_in_17_valid_a(array_11_io_d_in_17_valid_a),
    .io_d_in_17_b(array_11_io_d_in_17_b),
    .io_d_in_18_a(array_11_io_d_in_18_a),
    .io_d_in_18_valid_a(array_11_io_d_in_18_valid_a),
    .io_d_in_18_b(array_11_io_d_in_18_b),
    .io_d_in_19_a(array_11_io_d_in_19_a),
    .io_d_in_19_valid_a(array_11_io_d_in_19_valid_a),
    .io_d_in_19_b(array_11_io_d_in_19_b),
    .io_d_in_20_a(array_11_io_d_in_20_a),
    .io_d_in_20_valid_a(array_11_io_d_in_20_valid_a),
    .io_d_in_20_b(array_11_io_d_in_20_b),
    .io_d_in_21_a(array_11_io_d_in_21_a),
    .io_d_in_21_valid_a(array_11_io_d_in_21_valid_a),
    .io_d_in_21_b(array_11_io_d_in_21_b),
    .io_d_in_22_a(array_11_io_d_in_22_a),
    .io_d_in_22_valid_a(array_11_io_d_in_22_valid_a),
    .io_d_in_22_b(array_11_io_d_in_22_b),
    .io_d_in_23_a(array_11_io_d_in_23_a),
    .io_d_in_23_valid_a(array_11_io_d_in_23_valid_a),
    .io_d_in_23_b(array_11_io_d_in_23_b),
    .io_d_in_24_a(array_11_io_d_in_24_a),
    .io_d_in_24_valid_a(array_11_io_d_in_24_valid_a),
    .io_d_in_24_b(array_11_io_d_in_24_b),
    .io_d_in_25_a(array_11_io_d_in_25_a),
    .io_d_in_25_valid_a(array_11_io_d_in_25_valid_a),
    .io_d_in_25_b(array_11_io_d_in_25_b),
    .io_d_in_26_a(array_11_io_d_in_26_a),
    .io_d_in_26_valid_a(array_11_io_d_in_26_valid_a),
    .io_d_in_26_b(array_11_io_d_in_26_b),
    .io_d_in_27_a(array_11_io_d_in_27_a),
    .io_d_in_27_valid_a(array_11_io_d_in_27_valid_a),
    .io_d_in_27_b(array_11_io_d_in_27_b),
    .io_d_in_28_a(array_11_io_d_in_28_a),
    .io_d_in_28_valid_a(array_11_io_d_in_28_valid_a),
    .io_d_in_28_b(array_11_io_d_in_28_b),
    .io_d_in_29_a(array_11_io_d_in_29_a),
    .io_d_in_29_valid_a(array_11_io_d_in_29_valid_a),
    .io_d_in_29_b(array_11_io_d_in_29_b),
    .io_d_in_30_a(array_11_io_d_in_30_a),
    .io_d_in_30_valid_a(array_11_io_d_in_30_valid_a),
    .io_d_in_30_b(array_11_io_d_in_30_b),
    .io_d_in_31_a(array_11_io_d_in_31_a),
    .io_d_in_31_valid_a(array_11_io_d_in_31_valid_a),
    .io_d_in_31_b(array_11_io_d_in_31_b),
    .io_d_out_0_a(array_11_io_d_out_0_a),
    .io_d_out_0_valid_a(array_11_io_d_out_0_valid_a),
    .io_d_out_0_b(array_11_io_d_out_0_b),
    .io_d_out_0_valid_b(array_11_io_d_out_0_valid_b),
    .io_d_out_1_a(array_11_io_d_out_1_a),
    .io_d_out_1_valid_a(array_11_io_d_out_1_valid_a),
    .io_d_out_1_b(array_11_io_d_out_1_b),
    .io_d_out_1_valid_b(array_11_io_d_out_1_valid_b),
    .io_d_out_2_a(array_11_io_d_out_2_a),
    .io_d_out_2_valid_a(array_11_io_d_out_2_valid_a),
    .io_d_out_2_b(array_11_io_d_out_2_b),
    .io_d_out_2_valid_b(array_11_io_d_out_2_valid_b),
    .io_d_out_3_a(array_11_io_d_out_3_a),
    .io_d_out_3_valid_a(array_11_io_d_out_3_valid_a),
    .io_d_out_3_b(array_11_io_d_out_3_b),
    .io_d_out_3_valid_b(array_11_io_d_out_3_valid_b),
    .io_d_out_4_a(array_11_io_d_out_4_a),
    .io_d_out_4_valid_a(array_11_io_d_out_4_valid_a),
    .io_d_out_4_b(array_11_io_d_out_4_b),
    .io_d_out_4_valid_b(array_11_io_d_out_4_valid_b),
    .io_d_out_5_a(array_11_io_d_out_5_a),
    .io_d_out_5_valid_a(array_11_io_d_out_5_valid_a),
    .io_d_out_5_b(array_11_io_d_out_5_b),
    .io_d_out_5_valid_b(array_11_io_d_out_5_valid_b),
    .io_d_out_6_a(array_11_io_d_out_6_a),
    .io_d_out_6_valid_a(array_11_io_d_out_6_valid_a),
    .io_d_out_6_b(array_11_io_d_out_6_b),
    .io_d_out_6_valid_b(array_11_io_d_out_6_valid_b),
    .io_d_out_7_a(array_11_io_d_out_7_a),
    .io_d_out_7_valid_a(array_11_io_d_out_7_valid_a),
    .io_d_out_7_b(array_11_io_d_out_7_b),
    .io_d_out_7_valid_b(array_11_io_d_out_7_valid_b),
    .io_d_out_8_a(array_11_io_d_out_8_a),
    .io_d_out_8_valid_a(array_11_io_d_out_8_valid_a),
    .io_d_out_8_b(array_11_io_d_out_8_b),
    .io_d_out_8_valid_b(array_11_io_d_out_8_valid_b),
    .io_d_out_9_a(array_11_io_d_out_9_a),
    .io_d_out_9_valid_a(array_11_io_d_out_9_valid_a),
    .io_d_out_9_b(array_11_io_d_out_9_b),
    .io_d_out_9_valid_b(array_11_io_d_out_9_valid_b),
    .io_d_out_10_a(array_11_io_d_out_10_a),
    .io_d_out_10_valid_a(array_11_io_d_out_10_valid_a),
    .io_d_out_10_b(array_11_io_d_out_10_b),
    .io_d_out_10_valid_b(array_11_io_d_out_10_valid_b),
    .io_d_out_11_a(array_11_io_d_out_11_a),
    .io_d_out_11_valid_a(array_11_io_d_out_11_valid_a),
    .io_d_out_11_b(array_11_io_d_out_11_b),
    .io_d_out_11_valid_b(array_11_io_d_out_11_valid_b),
    .io_d_out_12_a(array_11_io_d_out_12_a),
    .io_d_out_12_valid_a(array_11_io_d_out_12_valid_a),
    .io_d_out_12_b(array_11_io_d_out_12_b),
    .io_d_out_12_valid_b(array_11_io_d_out_12_valid_b),
    .io_d_out_13_a(array_11_io_d_out_13_a),
    .io_d_out_13_valid_a(array_11_io_d_out_13_valid_a),
    .io_d_out_13_b(array_11_io_d_out_13_b),
    .io_d_out_13_valid_b(array_11_io_d_out_13_valid_b),
    .io_d_out_14_a(array_11_io_d_out_14_a),
    .io_d_out_14_valid_a(array_11_io_d_out_14_valid_a),
    .io_d_out_14_b(array_11_io_d_out_14_b),
    .io_d_out_14_valid_b(array_11_io_d_out_14_valid_b),
    .io_d_out_15_a(array_11_io_d_out_15_a),
    .io_d_out_15_valid_a(array_11_io_d_out_15_valid_a),
    .io_d_out_15_b(array_11_io_d_out_15_b),
    .io_d_out_15_valid_b(array_11_io_d_out_15_valid_b),
    .io_d_out_16_a(array_11_io_d_out_16_a),
    .io_d_out_16_valid_a(array_11_io_d_out_16_valid_a),
    .io_d_out_16_b(array_11_io_d_out_16_b),
    .io_d_out_16_valid_b(array_11_io_d_out_16_valid_b),
    .io_d_out_17_a(array_11_io_d_out_17_a),
    .io_d_out_17_valid_a(array_11_io_d_out_17_valid_a),
    .io_d_out_17_b(array_11_io_d_out_17_b),
    .io_d_out_17_valid_b(array_11_io_d_out_17_valid_b),
    .io_d_out_18_a(array_11_io_d_out_18_a),
    .io_d_out_18_valid_a(array_11_io_d_out_18_valid_a),
    .io_d_out_18_b(array_11_io_d_out_18_b),
    .io_d_out_18_valid_b(array_11_io_d_out_18_valid_b),
    .io_d_out_19_a(array_11_io_d_out_19_a),
    .io_d_out_19_valid_a(array_11_io_d_out_19_valid_a),
    .io_d_out_19_b(array_11_io_d_out_19_b),
    .io_d_out_19_valid_b(array_11_io_d_out_19_valid_b),
    .io_d_out_20_a(array_11_io_d_out_20_a),
    .io_d_out_20_valid_a(array_11_io_d_out_20_valid_a),
    .io_d_out_20_b(array_11_io_d_out_20_b),
    .io_d_out_20_valid_b(array_11_io_d_out_20_valid_b),
    .io_d_out_21_a(array_11_io_d_out_21_a),
    .io_d_out_21_valid_a(array_11_io_d_out_21_valid_a),
    .io_d_out_21_b(array_11_io_d_out_21_b),
    .io_d_out_21_valid_b(array_11_io_d_out_21_valid_b),
    .io_d_out_22_a(array_11_io_d_out_22_a),
    .io_d_out_22_valid_a(array_11_io_d_out_22_valid_a),
    .io_d_out_22_b(array_11_io_d_out_22_b),
    .io_d_out_22_valid_b(array_11_io_d_out_22_valid_b),
    .io_d_out_23_a(array_11_io_d_out_23_a),
    .io_d_out_23_valid_a(array_11_io_d_out_23_valid_a),
    .io_d_out_23_b(array_11_io_d_out_23_b),
    .io_d_out_23_valid_b(array_11_io_d_out_23_valid_b),
    .io_d_out_24_a(array_11_io_d_out_24_a),
    .io_d_out_24_valid_a(array_11_io_d_out_24_valid_a),
    .io_d_out_24_b(array_11_io_d_out_24_b),
    .io_d_out_24_valid_b(array_11_io_d_out_24_valid_b),
    .io_d_out_25_a(array_11_io_d_out_25_a),
    .io_d_out_25_valid_a(array_11_io_d_out_25_valid_a),
    .io_d_out_25_b(array_11_io_d_out_25_b),
    .io_d_out_25_valid_b(array_11_io_d_out_25_valid_b),
    .io_d_out_26_a(array_11_io_d_out_26_a),
    .io_d_out_26_valid_a(array_11_io_d_out_26_valid_a),
    .io_d_out_26_b(array_11_io_d_out_26_b),
    .io_d_out_26_valid_b(array_11_io_d_out_26_valid_b),
    .io_d_out_27_a(array_11_io_d_out_27_a),
    .io_d_out_27_valid_a(array_11_io_d_out_27_valid_a),
    .io_d_out_27_b(array_11_io_d_out_27_b),
    .io_d_out_27_valid_b(array_11_io_d_out_27_valid_b),
    .io_d_out_28_a(array_11_io_d_out_28_a),
    .io_d_out_28_valid_a(array_11_io_d_out_28_valid_a),
    .io_d_out_28_b(array_11_io_d_out_28_b),
    .io_d_out_28_valid_b(array_11_io_d_out_28_valid_b),
    .io_d_out_29_a(array_11_io_d_out_29_a),
    .io_d_out_29_valid_a(array_11_io_d_out_29_valid_a),
    .io_d_out_29_b(array_11_io_d_out_29_b),
    .io_d_out_29_valid_b(array_11_io_d_out_29_valid_b),
    .io_d_out_30_a(array_11_io_d_out_30_a),
    .io_d_out_30_valid_a(array_11_io_d_out_30_valid_a),
    .io_d_out_30_b(array_11_io_d_out_30_b),
    .io_d_out_30_valid_b(array_11_io_d_out_30_valid_b),
    .io_d_out_31_a(array_11_io_d_out_31_a),
    .io_d_out_31_valid_a(array_11_io_d_out_31_valid_a),
    .io_d_out_31_b(array_11_io_d_out_31_b),
    .io_d_out_31_valid_b(array_11_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_11_io_wr_en_mem1),
    .io_wr_en_mem2(array_11_io_wr_en_mem2),
    .io_wr_en_mem3(array_11_io_wr_en_mem3),
    .io_wr_en_mem4(array_11_io_wr_en_mem4),
    .io_wr_en_mem5(array_11_io_wr_en_mem5),
    .io_wr_en_mem6(array_11_io_wr_en_mem6),
    .io_wr_instr_mem1(array_11_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_11_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_11_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_11_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_11_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_11_io_wr_instr_mem6),
    .io_PC1_in(array_11_io_PC1_in),
    .io_PC6_out(array_11_io_PC6_out),
    .io_Addr_in(array_11_io_Addr_in),
    .io_Addr_out(array_11_io_Addr_out),
    .io_Tag_in_Tag(array_11_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_11_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_11_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_11_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_12 ( // @[Array.scala 41:54]
    .clock(array_12_clock),
    .reset(array_12_reset),
    .io_d_in_0_a(array_12_io_d_in_0_a),
    .io_d_in_0_valid_a(array_12_io_d_in_0_valid_a),
    .io_d_in_0_b(array_12_io_d_in_0_b),
    .io_d_in_1_a(array_12_io_d_in_1_a),
    .io_d_in_1_valid_a(array_12_io_d_in_1_valid_a),
    .io_d_in_1_b(array_12_io_d_in_1_b),
    .io_d_in_2_a(array_12_io_d_in_2_a),
    .io_d_in_2_valid_a(array_12_io_d_in_2_valid_a),
    .io_d_in_2_b(array_12_io_d_in_2_b),
    .io_d_in_3_a(array_12_io_d_in_3_a),
    .io_d_in_3_valid_a(array_12_io_d_in_3_valid_a),
    .io_d_in_3_b(array_12_io_d_in_3_b),
    .io_d_in_4_a(array_12_io_d_in_4_a),
    .io_d_in_4_valid_a(array_12_io_d_in_4_valid_a),
    .io_d_in_4_b(array_12_io_d_in_4_b),
    .io_d_in_5_a(array_12_io_d_in_5_a),
    .io_d_in_5_valid_a(array_12_io_d_in_5_valid_a),
    .io_d_in_5_b(array_12_io_d_in_5_b),
    .io_d_in_6_a(array_12_io_d_in_6_a),
    .io_d_in_6_valid_a(array_12_io_d_in_6_valid_a),
    .io_d_in_6_b(array_12_io_d_in_6_b),
    .io_d_in_7_a(array_12_io_d_in_7_a),
    .io_d_in_7_valid_a(array_12_io_d_in_7_valid_a),
    .io_d_in_7_b(array_12_io_d_in_7_b),
    .io_d_in_8_a(array_12_io_d_in_8_a),
    .io_d_in_8_valid_a(array_12_io_d_in_8_valid_a),
    .io_d_in_8_b(array_12_io_d_in_8_b),
    .io_d_in_9_a(array_12_io_d_in_9_a),
    .io_d_in_9_valid_a(array_12_io_d_in_9_valid_a),
    .io_d_in_9_b(array_12_io_d_in_9_b),
    .io_d_in_10_a(array_12_io_d_in_10_a),
    .io_d_in_10_valid_a(array_12_io_d_in_10_valid_a),
    .io_d_in_10_b(array_12_io_d_in_10_b),
    .io_d_in_11_a(array_12_io_d_in_11_a),
    .io_d_in_11_valid_a(array_12_io_d_in_11_valid_a),
    .io_d_in_11_b(array_12_io_d_in_11_b),
    .io_d_in_12_a(array_12_io_d_in_12_a),
    .io_d_in_12_valid_a(array_12_io_d_in_12_valid_a),
    .io_d_in_12_b(array_12_io_d_in_12_b),
    .io_d_in_13_a(array_12_io_d_in_13_a),
    .io_d_in_13_valid_a(array_12_io_d_in_13_valid_a),
    .io_d_in_13_b(array_12_io_d_in_13_b),
    .io_d_in_14_a(array_12_io_d_in_14_a),
    .io_d_in_14_valid_a(array_12_io_d_in_14_valid_a),
    .io_d_in_14_b(array_12_io_d_in_14_b),
    .io_d_in_15_a(array_12_io_d_in_15_a),
    .io_d_in_15_valid_a(array_12_io_d_in_15_valid_a),
    .io_d_in_15_b(array_12_io_d_in_15_b),
    .io_d_in_16_a(array_12_io_d_in_16_a),
    .io_d_in_16_valid_a(array_12_io_d_in_16_valid_a),
    .io_d_in_16_b(array_12_io_d_in_16_b),
    .io_d_in_17_a(array_12_io_d_in_17_a),
    .io_d_in_17_valid_a(array_12_io_d_in_17_valid_a),
    .io_d_in_17_b(array_12_io_d_in_17_b),
    .io_d_in_18_a(array_12_io_d_in_18_a),
    .io_d_in_18_valid_a(array_12_io_d_in_18_valid_a),
    .io_d_in_18_b(array_12_io_d_in_18_b),
    .io_d_in_19_a(array_12_io_d_in_19_a),
    .io_d_in_19_valid_a(array_12_io_d_in_19_valid_a),
    .io_d_in_19_b(array_12_io_d_in_19_b),
    .io_d_in_20_a(array_12_io_d_in_20_a),
    .io_d_in_20_valid_a(array_12_io_d_in_20_valid_a),
    .io_d_in_20_b(array_12_io_d_in_20_b),
    .io_d_in_21_a(array_12_io_d_in_21_a),
    .io_d_in_21_valid_a(array_12_io_d_in_21_valid_a),
    .io_d_in_21_b(array_12_io_d_in_21_b),
    .io_d_in_22_a(array_12_io_d_in_22_a),
    .io_d_in_22_valid_a(array_12_io_d_in_22_valid_a),
    .io_d_in_22_b(array_12_io_d_in_22_b),
    .io_d_in_23_a(array_12_io_d_in_23_a),
    .io_d_in_23_valid_a(array_12_io_d_in_23_valid_a),
    .io_d_in_23_b(array_12_io_d_in_23_b),
    .io_d_in_24_a(array_12_io_d_in_24_a),
    .io_d_in_24_valid_a(array_12_io_d_in_24_valid_a),
    .io_d_in_24_b(array_12_io_d_in_24_b),
    .io_d_in_25_a(array_12_io_d_in_25_a),
    .io_d_in_25_valid_a(array_12_io_d_in_25_valid_a),
    .io_d_in_25_b(array_12_io_d_in_25_b),
    .io_d_in_26_a(array_12_io_d_in_26_a),
    .io_d_in_26_valid_a(array_12_io_d_in_26_valid_a),
    .io_d_in_26_b(array_12_io_d_in_26_b),
    .io_d_in_27_a(array_12_io_d_in_27_a),
    .io_d_in_27_valid_a(array_12_io_d_in_27_valid_a),
    .io_d_in_27_b(array_12_io_d_in_27_b),
    .io_d_in_28_a(array_12_io_d_in_28_a),
    .io_d_in_28_valid_a(array_12_io_d_in_28_valid_a),
    .io_d_in_28_b(array_12_io_d_in_28_b),
    .io_d_in_29_a(array_12_io_d_in_29_a),
    .io_d_in_29_valid_a(array_12_io_d_in_29_valid_a),
    .io_d_in_29_b(array_12_io_d_in_29_b),
    .io_d_in_30_a(array_12_io_d_in_30_a),
    .io_d_in_30_valid_a(array_12_io_d_in_30_valid_a),
    .io_d_in_30_b(array_12_io_d_in_30_b),
    .io_d_in_31_a(array_12_io_d_in_31_a),
    .io_d_in_31_valid_a(array_12_io_d_in_31_valid_a),
    .io_d_in_31_b(array_12_io_d_in_31_b),
    .io_d_out_0_a(array_12_io_d_out_0_a),
    .io_d_out_0_valid_a(array_12_io_d_out_0_valid_a),
    .io_d_out_0_b(array_12_io_d_out_0_b),
    .io_d_out_0_valid_b(array_12_io_d_out_0_valid_b),
    .io_d_out_1_a(array_12_io_d_out_1_a),
    .io_d_out_1_valid_a(array_12_io_d_out_1_valid_a),
    .io_d_out_1_b(array_12_io_d_out_1_b),
    .io_d_out_1_valid_b(array_12_io_d_out_1_valid_b),
    .io_d_out_2_a(array_12_io_d_out_2_a),
    .io_d_out_2_valid_a(array_12_io_d_out_2_valid_a),
    .io_d_out_2_b(array_12_io_d_out_2_b),
    .io_d_out_2_valid_b(array_12_io_d_out_2_valid_b),
    .io_d_out_3_a(array_12_io_d_out_3_a),
    .io_d_out_3_valid_a(array_12_io_d_out_3_valid_a),
    .io_d_out_3_b(array_12_io_d_out_3_b),
    .io_d_out_3_valid_b(array_12_io_d_out_3_valid_b),
    .io_d_out_4_a(array_12_io_d_out_4_a),
    .io_d_out_4_valid_a(array_12_io_d_out_4_valid_a),
    .io_d_out_4_b(array_12_io_d_out_4_b),
    .io_d_out_4_valid_b(array_12_io_d_out_4_valid_b),
    .io_d_out_5_a(array_12_io_d_out_5_a),
    .io_d_out_5_valid_a(array_12_io_d_out_5_valid_a),
    .io_d_out_5_b(array_12_io_d_out_5_b),
    .io_d_out_5_valid_b(array_12_io_d_out_5_valid_b),
    .io_d_out_6_a(array_12_io_d_out_6_a),
    .io_d_out_6_valid_a(array_12_io_d_out_6_valid_a),
    .io_d_out_6_b(array_12_io_d_out_6_b),
    .io_d_out_6_valid_b(array_12_io_d_out_6_valid_b),
    .io_d_out_7_a(array_12_io_d_out_7_a),
    .io_d_out_7_valid_a(array_12_io_d_out_7_valid_a),
    .io_d_out_7_b(array_12_io_d_out_7_b),
    .io_d_out_7_valid_b(array_12_io_d_out_7_valid_b),
    .io_d_out_8_a(array_12_io_d_out_8_a),
    .io_d_out_8_valid_a(array_12_io_d_out_8_valid_a),
    .io_d_out_8_b(array_12_io_d_out_8_b),
    .io_d_out_8_valid_b(array_12_io_d_out_8_valid_b),
    .io_d_out_9_a(array_12_io_d_out_9_a),
    .io_d_out_9_valid_a(array_12_io_d_out_9_valid_a),
    .io_d_out_9_b(array_12_io_d_out_9_b),
    .io_d_out_9_valid_b(array_12_io_d_out_9_valid_b),
    .io_d_out_10_a(array_12_io_d_out_10_a),
    .io_d_out_10_valid_a(array_12_io_d_out_10_valid_a),
    .io_d_out_10_b(array_12_io_d_out_10_b),
    .io_d_out_10_valid_b(array_12_io_d_out_10_valid_b),
    .io_d_out_11_a(array_12_io_d_out_11_a),
    .io_d_out_11_valid_a(array_12_io_d_out_11_valid_a),
    .io_d_out_11_b(array_12_io_d_out_11_b),
    .io_d_out_11_valid_b(array_12_io_d_out_11_valid_b),
    .io_d_out_12_a(array_12_io_d_out_12_a),
    .io_d_out_12_valid_a(array_12_io_d_out_12_valid_a),
    .io_d_out_12_b(array_12_io_d_out_12_b),
    .io_d_out_12_valid_b(array_12_io_d_out_12_valid_b),
    .io_d_out_13_a(array_12_io_d_out_13_a),
    .io_d_out_13_valid_a(array_12_io_d_out_13_valid_a),
    .io_d_out_13_b(array_12_io_d_out_13_b),
    .io_d_out_13_valid_b(array_12_io_d_out_13_valid_b),
    .io_d_out_14_a(array_12_io_d_out_14_a),
    .io_d_out_14_valid_a(array_12_io_d_out_14_valid_a),
    .io_d_out_14_b(array_12_io_d_out_14_b),
    .io_d_out_14_valid_b(array_12_io_d_out_14_valid_b),
    .io_d_out_15_a(array_12_io_d_out_15_a),
    .io_d_out_15_valid_a(array_12_io_d_out_15_valid_a),
    .io_d_out_15_b(array_12_io_d_out_15_b),
    .io_d_out_15_valid_b(array_12_io_d_out_15_valid_b),
    .io_d_out_16_a(array_12_io_d_out_16_a),
    .io_d_out_16_valid_a(array_12_io_d_out_16_valid_a),
    .io_d_out_16_b(array_12_io_d_out_16_b),
    .io_d_out_16_valid_b(array_12_io_d_out_16_valid_b),
    .io_d_out_17_a(array_12_io_d_out_17_a),
    .io_d_out_17_valid_a(array_12_io_d_out_17_valid_a),
    .io_d_out_17_b(array_12_io_d_out_17_b),
    .io_d_out_17_valid_b(array_12_io_d_out_17_valid_b),
    .io_d_out_18_a(array_12_io_d_out_18_a),
    .io_d_out_18_valid_a(array_12_io_d_out_18_valid_a),
    .io_d_out_18_b(array_12_io_d_out_18_b),
    .io_d_out_18_valid_b(array_12_io_d_out_18_valid_b),
    .io_d_out_19_a(array_12_io_d_out_19_a),
    .io_d_out_19_valid_a(array_12_io_d_out_19_valid_a),
    .io_d_out_19_b(array_12_io_d_out_19_b),
    .io_d_out_19_valid_b(array_12_io_d_out_19_valid_b),
    .io_d_out_20_a(array_12_io_d_out_20_a),
    .io_d_out_20_valid_a(array_12_io_d_out_20_valid_a),
    .io_d_out_20_b(array_12_io_d_out_20_b),
    .io_d_out_20_valid_b(array_12_io_d_out_20_valid_b),
    .io_d_out_21_a(array_12_io_d_out_21_a),
    .io_d_out_21_valid_a(array_12_io_d_out_21_valid_a),
    .io_d_out_21_b(array_12_io_d_out_21_b),
    .io_d_out_21_valid_b(array_12_io_d_out_21_valid_b),
    .io_d_out_22_a(array_12_io_d_out_22_a),
    .io_d_out_22_valid_a(array_12_io_d_out_22_valid_a),
    .io_d_out_22_b(array_12_io_d_out_22_b),
    .io_d_out_22_valid_b(array_12_io_d_out_22_valid_b),
    .io_d_out_23_a(array_12_io_d_out_23_a),
    .io_d_out_23_valid_a(array_12_io_d_out_23_valid_a),
    .io_d_out_23_b(array_12_io_d_out_23_b),
    .io_d_out_23_valid_b(array_12_io_d_out_23_valid_b),
    .io_d_out_24_a(array_12_io_d_out_24_a),
    .io_d_out_24_valid_a(array_12_io_d_out_24_valid_a),
    .io_d_out_24_b(array_12_io_d_out_24_b),
    .io_d_out_24_valid_b(array_12_io_d_out_24_valid_b),
    .io_d_out_25_a(array_12_io_d_out_25_a),
    .io_d_out_25_valid_a(array_12_io_d_out_25_valid_a),
    .io_d_out_25_b(array_12_io_d_out_25_b),
    .io_d_out_25_valid_b(array_12_io_d_out_25_valid_b),
    .io_d_out_26_a(array_12_io_d_out_26_a),
    .io_d_out_26_valid_a(array_12_io_d_out_26_valid_a),
    .io_d_out_26_b(array_12_io_d_out_26_b),
    .io_d_out_26_valid_b(array_12_io_d_out_26_valid_b),
    .io_d_out_27_a(array_12_io_d_out_27_a),
    .io_d_out_27_valid_a(array_12_io_d_out_27_valid_a),
    .io_d_out_27_b(array_12_io_d_out_27_b),
    .io_d_out_27_valid_b(array_12_io_d_out_27_valid_b),
    .io_d_out_28_a(array_12_io_d_out_28_a),
    .io_d_out_28_valid_a(array_12_io_d_out_28_valid_a),
    .io_d_out_28_b(array_12_io_d_out_28_b),
    .io_d_out_28_valid_b(array_12_io_d_out_28_valid_b),
    .io_d_out_29_a(array_12_io_d_out_29_a),
    .io_d_out_29_valid_a(array_12_io_d_out_29_valid_a),
    .io_d_out_29_b(array_12_io_d_out_29_b),
    .io_d_out_29_valid_b(array_12_io_d_out_29_valid_b),
    .io_d_out_30_a(array_12_io_d_out_30_a),
    .io_d_out_30_valid_a(array_12_io_d_out_30_valid_a),
    .io_d_out_30_b(array_12_io_d_out_30_b),
    .io_d_out_30_valid_b(array_12_io_d_out_30_valid_b),
    .io_d_out_31_a(array_12_io_d_out_31_a),
    .io_d_out_31_valid_a(array_12_io_d_out_31_valid_a),
    .io_d_out_31_b(array_12_io_d_out_31_b),
    .io_d_out_31_valid_b(array_12_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_12_io_wr_en_mem1),
    .io_wr_en_mem2(array_12_io_wr_en_mem2),
    .io_wr_en_mem3(array_12_io_wr_en_mem3),
    .io_wr_en_mem4(array_12_io_wr_en_mem4),
    .io_wr_en_mem5(array_12_io_wr_en_mem5),
    .io_wr_en_mem6(array_12_io_wr_en_mem6),
    .io_wr_instr_mem1(array_12_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_12_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_12_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_12_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_12_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_12_io_wr_instr_mem6),
    .io_PC1_in(array_12_io_PC1_in),
    .io_PC6_out(array_12_io_PC6_out),
    .io_Addr_in(array_12_io_Addr_in),
    .io_Addr_out(array_12_io_Addr_out),
    .io_Tag_in_Tag(array_12_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_12_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_12_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_12_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_13 ( // @[Array.scala 41:54]
    .clock(array_13_clock),
    .reset(array_13_reset),
    .io_d_in_0_a(array_13_io_d_in_0_a),
    .io_d_in_0_valid_a(array_13_io_d_in_0_valid_a),
    .io_d_in_0_b(array_13_io_d_in_0_b),
    .io_d_in_1_a(array_13_io_d_in_1_a),
    .io_d_in_1_valid_a(array_13_io_d_in_1_valid_a),
    .io_d_in_1_b(array_13_io_d_in_1_b),
    .io_d_in_2_a(array_13_io_d_in_2_a),
    .io_d_in_2_valid_a(array_13_io_d_in_2_valid_a),
    .io_d_in_2_b(array_13_io_d_in_2_b),
    .io_d_in_3_a(array_13_io_d_in_3_a),
    .io_d_in_3_valid_a(array_13_io_d_in_3_valid_a),
    .io_d_in_3_b(array_13_io_d_in_3_b),
    .io_d_in_4_a(array_13_io_d_in_4_a),
    .io_d_in_4_valid_a(array_13_io_d_in_4_valid_a),
    .io_d_in_4_b(array_13_io_d_in_4_b),
    .io_d_in_5_a(array_13_io_d_in_5_a),
    .io_d_in_5_valid_a(array_13_io_d_in_5_valid_a),
    .io_d_in_5_b(array_13_io_d_in_5_b),
    .io_d_in_6_a(array_13_io_d_in_6_a),
    .io_d_in_6_valid_a(array_13_io_d_in_6_valid_a),
    .io_d_in_6_b(array_13_io_d_in_6_b),
    .io_d_in_7_a(array_13_io_d_in_7_a),
    .io_d_in_7_valid_a(array_13_io_d_in_7_valid_a),
    .io_d_in_7_b(array_13_io_d_in_7_b),
    .io_d_in_8_a(array_13_io_d_in_8_a),
    .io_d_in_8_valid_a(array_13_io_d_in_8_valid_a),
    .io_d_in_8_b(array_13_io_d_in_8_b),
    .io_d_in_9_a(array_13_io_d_in_9_a),
    .io_d_in_9_valid_a(array_13_io_d_in_9_valid_a),
    .io_d_in_9_b(array_13_io_d_in_9_b),
    .io_d_in_10_a(array_13_io_d_in_10_a),
    .io_d_in_10_valid_a(array_13_io_d_in_10_valid_a),
    .io_d_in_10_b(array_13_io_d_in_10_b),
    .io_d_in_11_a(array_13_io_d_in_11_a),
    .io_d_in_11_valid_a(array_13_io_d_in_11_valid_a),
    .io_d_in_11_b(array_13_io_d_in_11_b),
    .io_d_in_12_a(array_13_io_d_in_12_a),
    .io_d_in_12_valid_a(array_13_io_d_in_12_valid_a),
    .io_d_in_12_b(array_13_io_d_in_12_b),
    .io_d_in_13_a(array_13_io_d_in_13_a),
    .io_d_in_13_valid_a(array_13_io_d_in_13_valid_a),
    .io_d_in_13_b(array_13_io_d_in_13_b),
    .io_d_in_14_a(array_13_io_d_in_14_a),
    .io_d_in_14_valid_a(array_13_io_d_in_14_valid_a),
    .io_d_in_14_b(array_13_io_d_in_14_b),
    .io_d_in_15_a(array_13_io_d_in_15_a),
    .io_d_in_15_valid_a(array_13_io_d_in_15_valid_a),
    .io_d_in_15_b(array_13_io_d_in_15_b),
    .io_d_in_16_a(array_13_io_d_in_16_a),
    .io_d_in_16_valid_a(array_13_io_d_in_16_valid_a),
    .io_d_in_16_b(array_13_io_d_in_16_b),
    .io_d_in_17_a(array_13_io_d_in_17_a),
    .io_d_in_17_valid_a(array_13_io_d_in_17_valid_a),
    .io_d_in_17_b(array_13_io_d_in_17_b),
    .io_d_in_18_a(array_13_io_d_in_18_a),
    .io_d_in_18_valid_a(array_13_io_d_in_18_valid_a),
    .io_d_in_18_b(array_13_io_d_in_18_b),
    .io_d_in_19_a(array_13_io_d_in_19_a),
    .io_d_in_19_valid_a(array_13_io_d_in_19_valid_a),
    .io_d_in_19_b(array_13_io_d_in_19_b),
    .io_d_in_20_a(array_13_io_d_in_20_a),
    .io_d_in_20_valid_a(array_13_io_d_in_20_valid_a),
    .io_d_in_20_b(array_13_io_d_in_20_b),
    .io_d_in_21_a(array_13_io_d_in_21_a),
    .io_d_in_21_valid_a(array_13_io_d_in_21_valid_a),
    .io_d_in_21_b(array_13_io_d_in_21_b),
    .io_d_in_22_a(array_13_io_d_in_22_a),
    .io_d_in_22_valid_a(array_13_io_d_in_22_valid_a),
    .io_d_in_22_b(array_13_io_d_in_22_b),
    .io_d_in_23_a(array_13_io_d_in_23_a),
    .io_d_in_23_valid_a(array_13_io_d_in_23_valid_a),
    .io_d_in_23_b(array_13_io_d_in_23_b),
    .io_d_in_24_a(array_13_io_d_in_24_a),
    .io_d_in_24_valid_a(array_13_io_d_in_24_valid_a),
    .io_d_in_24_b(array_13_io_d_in_24_b),
    .io_d_in_25_a(array_13_io_d_in_25_a),
    .io_d_in_25_valid_a(array_13_io_d_in_25_valid_a),
    .io_d_in_25_b(array_13_io_d_in_25_b),
    .io_d_in_26_a(array_13_io_d_in_26_a),
    .io_d_in_26_valid_a(array_13_io_d_in_26_valid_a),
    .io_d_in_26_b(array_13_io_d_in_26_b),
    .io_d_in_27_a(array_13_io_d_in_27_a),
    .io_d_in_27_valid_a(array_13_io_d_in_27_valid_a),
    .io_d_in_27_b(array_13_io_d_in_27_b),
    .io_d_in_28_a(array_13_io_d_in_28_a),
    .io_d_in_28_valid_a(array_13_io_d_in_28_valid_a),
    .io_d_in_28_b(array_13_io_d_in_28_b),
    .io_d_in_29_a(array_13_io_d_in_29_a),
    .io_d_in_29_valid_a(array_13_io_d_in_29_valid_a),
    .io_d_in_29_b(array_13_io_d_in_29_b),
    .io_d_in_30_a(array_13_io_d_in_30_a),
    .io_d_in_30_valid_a(array_13_io_d_in_30_valid_a),
    .io_d_in_30_b(array_13_io_d_in_30_b),
    .io_d_in_31_a(array_13_io_d_in_31_a),
    .io_d_in_31_valid_a(array_13_io_d_in_31_valid_a),
    .io_d_in_31_b(array_13_io_d_in_31_b),
    .io_d_out_0_a(array_13_io_d_out_0_a),
    .io_d_out_0_valid_a(array_13_io_d_out_0_valid_a),
    .io_d_out_0_b(array_13_io_d_out_0_b),
    .io_d_out_0_valid_b(array_13_io_d_out_0_valid_b),
    .io_d_out_1_a(array_13_io_d_out_1_a),
    .io_d_out_1_valid_a(array_13_io_d_out_1_valid_a),
    .io_d_out_1_b(array_13_io_d_out_1_b),
    .io_d_out_1_valid_b(array_13_io_d_out_1_valid_b),
    .io_d_out_2_a(array_13_io_d_out_2_a),
    .io_d_out_2_valid_a(array_13_io_d_out_2_valid_a),
    .io_d_out_2_b(array_13_io_d_out_2_b),
    .io_d_out_2_valid_b(array_13_io_d_out_2_valid_b),
    .io_d_out_3_a(array_13_io_d_out_3_a),
    .io_d_out_3_valid_a(array_13_io_d_out_3_valid_a),
    .io_d_out_3_b(array_13_io_d_out_3_b),
    .io_d_out_3_valid_b(array_13_io_d_out_3_valid_b),
    .io_d_out_4_a(array_13_io_d_out_4_a),
    .io_d_out_4_valid_a(array_13_io_d_out_4_valid_a),
    .io_d_out_4_b(array_13_io_d_out_4_b),
    .io_d_out_4_valid_b(array_13_io_d_out_4_valid_b),
    .io_d_out_5_a(array_13_io_d_out_5_a),
    .io_d_out_5_valid_a(array_13_io_d_out_5_valid_a),
    .io_d_out_5_b(array_13_io_d_out_5_b),
    .io_d_out_5_valid_b(array_13_io_d_out_5_valid_b),
    .io_d_out_6_a(array_13_io_d_out_6_a),
    .io_d_out_6_valid_a(array_13_io_d_out_6_valid_a),
    .io_d_out_6_b(array_13_io_d_out_6_b),
    .io_d_out_6_valid_b(array_13_io_d_out_6_valid_b),
    .io_d_out_7_a(array_13_io_d_out_7_a),
    .io_d_out_7_valid_a(array_13_io_d_out_7_valid_a),
    .io_d_out_7_b(array_13_io_d_out_7_b),
    .io_d_out_7_valid_b(array_13_io_d_out_7_valid_b),
    .io_d_out_8_a(array_13_io_d_out_8_a),
    .io_d_out_8_valid_a(array_13_io_d_out_8_valid_a),
    .io_d_out_8_b(array_13_io_d_out_8_b),
    .io_d_out_8_valid_b(array_13_io_d_out_8_valid_b),
    .io_d_out_9_a(array_13_io_d_out_9_a),
    .io_d_out_9_valid_a(array_13_io_d_out_9_valid_a),
    .io_d_out_9_b(array_13_io_d_out_9_b),
    .io_d_out_9_valid_b(array_13_io_d_out_9_valid_b),
    .io_d_out_10_a(array_13_io_d_out_10_a),
    .io_d_out_10_valid_a(array_13_io_d_out_10_valid_a),
    .io_d_out_10_b(array_13_io_d_out_10_b),
    .io_d_out_10_valid_b(array_13_io_d_out_10_valid_b),
    .io_d_out_11_a(array_13_io_d_out_11_a),
    .io_d_out_11_valid_a(array_13_io_d_out_11_valid_a),
    .io_d_out_11_b(array_13_io_d_out_11_b),
    .io_d_out_11_valid_b(array_13_io_d_out_11_valid_b),
    .io_d_out_12_a(array_13_io_d_out_12_a),
    .io_d_out_12_valid_a(array_13_io_d_out_12_valid_a),
    .io_d_out_12_b(array_13_io_d_out_12_b),
    .io_d_out_12_valid_b(array_13_io_d_out_12_valid_b),
    .io_d_out_13_a(array_13_io_d_out_13_a),
    .io_d_out_13_valid_a(array_13_io_d_out_13_valid_a),
    .io_d_out_13_b(array_13_io_d_out_13_b),
    .io_d_out_13_valid_b(array_13_io_d_out_13_valid_b),
    .io_d_out_14_a(array_13_io_d_out_14_a),
    .io_d_out_14_valid_a(array_13_io_d_out_14_valid_a),
    .io_d_out_14_b(array_13_io_d_out_14_b),
    .io_d_out_14_valid_b(array_13_io_d_out_14_valid_b),
    .io_d_out_15_a(array_13_io_d_out_15_a),
    .io_d_out_15_valid_a(array_13_io_d_out_15_valid_a),
    .io_d_out_15_b(array_13_io_d_out_15_b),
    .io_d_out_15_valid_b(array_13_io_d_out_15_valid_b),
    .io_d_out_16_a(array_13_io_d_out_16_a),
    .io_d_out_16_valid_a(array_13_io_d_out_16_valid_a),
    .io_d_out_16_b(array_13_io_d_out_16_b),
    .io_d_out_16_valid_b(array_13_io_d_out_16_valid_b),
    .io_d_out_17_a(array_13_io_d_out_17_a),
    .io_d_out_17_valid_a(array_13_io_d_out_17_valid_a),
    .io_d_out_17_b(array_13_io_d_out_17_b),
    .io_d_out_17_valid_b(array_13_io_d_out_17_valid_b),
    .io_d_out_18_a(array_13_io_d_out_18_a),
    .io_d_out_18_valid_a(array_13_io_d_out_18_valid_a),
    .io_d_out_18_b(array_13_io_d_out_18_b),
    .io_d_out_18_valid_b(array_13_io_d_out_18_valid_b),
    .io_d_out_19_a(array_13_io_d_out_19_a),
    .io_d_out_19_valid_a(array_13_io_d_out_19_valid_a),
    .io_d_out_19_b(array_13_io_d_out_19_b),
    .io_d_out_19_valid_b(array_13_io_d_out_19_valid_b),
    .io_d_out_20_a(array_13_io_d_out_20_a),
    .io_d_out_20_valid_a(array_13_io_d_out_20_valid_a),
    .io_d_out_20_b(array_13_io_d_out_20_b),
    .io_d_out_20_valid_b(array_13_io_d_out_20_valid_b),
    .io_d_out_21_a(array_13_io_d_out_21_a),
    .io_d_out_21_valid_a(array_13_io_d_out_21_valid_a),
    .io_d_out_21_b(array_13_io_d_out_21_b),
    .io_d_out_21_valid_b(array_13_io_d_out_21_valid_b),
    .io_d_out_22_a(array_13_io_d_out_22_a),
    .io_d_out_22_valid_a(array_13_io_d_out_22_valid_a),
    .io_d_out_22_b(array_13_io_d_out_22_b),
    .io_d_out_22_valid_b(array_13_io_d_out_22_valid_b),
    .io_d_out_23_a(array_13_io_d_out_23_a),
    .io_d_out_23_valid_a(array_13_io_d_out_23_valid_a),
    .io_d_out_23_b(array_13_io_d_out_23_b),
    .io_d_out_23_valid_b(array_13_io_d_out_23_valid_b),
    .io_d_out_24_a(array_13_io_d_out_24_a),
    .io_d_out_24_valid_a(array_13_io_d_out_24_valid_a),
    .io_d_out_24_b(array_13_io_d_out_24_b),
    .io_d_out_24_valid_b(array_13_io_d_out_24_valid_b),
    .io_d_out_25_a(array_13_io_d_out_25_a),
    .io_d_out_25_valid_a(array_13_io_d_out_25_valid_a),
    .io_d_out_25_b(array_13_io_d_out_25_b),
    .io_d_out_25_valid_b(array_13_io_d_out_25_valid_b),
    .io_d_out_26_a(array_13_io_d_out_26_a),
    .io_d_out_26_valid_a(array_13_io_d_out_26_valid_a),
    .io_d_out_26_b(array_13_io_d_out_26_b),
    .io_d_out_26_valid_b(array_13_io_d_out_26_valid_b),
    .io_d_out_27_a(array_13_io_d_out_27_a),
    .io_d_out_27_valid_a(array_13_io_d_out_27_valid_a),
    .io_d_out_27_b(array_13_io_d_out_27_b),
    .io_d_out_27_valid_b(array_13_io_d_out_27_valid_b),
    .io_d_out_28_a(array_13_io_d_out_28_a),
    .io_d_out_28_valid_a(array_13_io_d_out_28_valid_a),
    .io_d_out_28_b(array_13_io_d_out_28_b),
    .io_d_out_28_valid_b(array_13_io_d_out_28_valid_b),
    .io_d_out_29_a(array_13_io_d_out_29_a),
    .io_d_out_29_valid_a(array_13_io_d_out_29_valid_a),
    .io_d_out_29_b(array_13_io_d_out_29_b),
    .io_d_out_29_valid_b(array_13_io_d_out_29_valid_b),
    .io_d_out_30_a(array_13_io_d_out_30_a),
    .io_d_out_30_valid_a(array_13_io_d_out_30_valid_a),
    .io_d_out_30_b(array_13_io_d_out_30_b),
    .io_d_out_30_valid_b(array_13_io_d_out_30_valid_b),
    .io_d_out_31_a(array_13_io_d_out_31_a),
    .io_d_out_31_valid_a(array_13_io_d_out_31_valid_a),
    .io_d_out_31_b(array_13_io_d_out_31_b),
    .io_d_out_31_valid_b(array_13_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_13_io_wr_en_mem1),
    .io_wr_en_mem2(array_13_io_wr_en_mem2),
    .io_wr_en_mem3(array_13_io_wr_en_mem3),
    .io_wr_en_mem4(array_13_io_wr_en_mem4),
    .io_wr_en_mem5(array_13_io_wr_en_mem5),
    .io_wr_en_mem6(array_13_io_wr_en_mem6),
    .io_wr_instr_mem1(array_13_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_13_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_13_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_13_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_13_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_13_io_wr_instr_mem6),
    .io_PC1_in(array_13_io_PC1_in),
    .io_PC6_out(array_13_io_PC6_out),
    .io_Addr_in(array_13_io_Addr_in),
    .io_Addr_out(array_13_io_Addr_out),
    .io_Tag_in_Tag(array_13_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_13_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_13_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_13_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_14 ( // @[Array.scala 41:54]
    .clock(array_14_clock),
    .reset(array_14_reset),
    .io_d_in_0_a(array_14_io_d_in_0_a),
    .io_d_in_0_valid_a(array_14_io_d_in_0_valid_a),
    .io_d_in_0_b(array_14_io_d_in_0_b),
    .io_d_in_1_a(array_14_io_d_in_1_a),
    .io_d_in_1_valid_a(array_14_io_d_in_1_valid_a),
    .io_d_in_1_b(array_14_io_d_in_1_b),
    .io_d_in_2_a(array_14_io_d_in_2_a),
    .io_d_in_2_valid_a(array_14_io_d_in_2_valid_a),
    .io_d_in_2_b(array_14_io_d_in_2_b),
    .io_d_in_3_a(array_14_io_d_in_3_a),
    .io_d_in_3_valid_a(array_14_io_d_in_3_valid_a),
    .io_d_in_3_b(array_14_io_d_in_3_b),
    .io_d_in_4_a(array_14_io_d_in_4_a),
    .io_d_in_4_valid_a(array_14_io_d_in_4_valid_a),
    .io_d_in_4_b(array_14_io_d_in_4_b),
    .io_d_in_5_a(array_14_io_d_in_5_a),
    .io_d_in_5_valid_a(array_14_io_d_in_5_valid_a),
    .io_d_in_5_b(array_14_io_d_in_5_b),
    .io_d_in_6_a(array_14_io_d_in_6_a),
    .io_d_in_6_valid_a(array_14_io_d_in_6_valid_a),
    .io_d_in_6_b(array_14_io_d_in_6_b),
    .io_d_in_7_a(array_14_io_d_in_7_a),
    .io_d_in_7_valid_a(array_14_io_d_in_7_valid_a),
    .io_d_in_7_b(array_14_io_d_in_7_b),
    .io_d_in_8_a(array_14_io_d_in_8_a),
    .io_d_in_8_valid_a(array_14_io_d_in_8_valid_a),
    .io_d_in_8_b(array_14_io_d_in_8_b),
    .io_d_in_9_a(array_14_io_d_in_9_a),
    .io_d_in_9_valid_a(array_14_io_d_in_9_valid_a),
    .io_d_in_9_b(array_14_io_d_in_9_b),
    .io_d_in_10_a(array_14_io_d_in_10_a),
    .io_d_in_10_valid_a(array_14_io_d_in_10_valid_a),
    .io_d_in_10_b(array_14_io_d_in_10_b),
    .io_d_in_11_a(array_14_io_d_in_11_a),
    .io_d_in_11_valid_a(array_14_io_d_in_11_valid_a),
    .io_d_in_11_b(array_14_io_d_in_11_b),
    .io_d_in_12_a(array_14_io_d_in_12_a),
    .io_d_in_12_valid_a(array_14_io_d_in_12_valid_a),
    .io_d_in_12_b(array_14_io_d_in_12_b),
    .io_d_in_13_a(array_14_io_d_in_13_a),
    .io_d_in_13_valid_a(array_14_io_d_in_13_valid_a),
    .io_d_in_13_b(array_14_io_d_in_13_b),
    .io_d_in_14_a(array_14_io_d_in_14_a),
    .io_d_in_14_valid_a(array_14_io_d_in_14_valid_a),
    .io_d_in_14_b(array_14_io_d_in_14_b),
    .io_d_in_15_a(array_14_io_d_in_15_a),
    .io_d_in_15_valid_a(array_14_io_d_in_15_valid_a),
    .io_d_in_15_b(array_14_io_d_in_15_b),
    .io_d_in_16_a(array_14_io_d_in_16_a),
    .io_d_in_16_valid_a(array_14_io_d_in_16_valid_a),
    .io_d_in_16_b(array_14_io_d_in_16_b),
    .io_d_in_17_a(array_14_io_d_in_17_a),
    .io_d_in_17_valid_a(array_14_io_d_in_17_valid_a),
    .io_d_in_17_b(array_14_io_d_in_17_b),
    .io_d_in_18_a(array_14_io_d_in_18_a),
    .io_d_in_18_valid_a(array_14_io_d_in_18_valid_a),
    .io_d_in_18_b(array_14_io_d_in_18_b),
    .io_d_in_19_a(array_14_io_d_in_19_a),
    .io_d_in_19_valid_a(array_14_io_d_in_19_valid_a),
    .io_d_in_19_b(array_14_io_d_in_19_b),
    .io_d_in_20_a(array_14_io_d_in_20_a),
    .io_d_in_20_valid_a(array_14_io_d_in_20_valid_a),
    .io_d_in_20_b(array_14_io_d_in_20_b),
    .io_d_in_21_a(array_14_io_d_in_21_a),
    .io_d_in_21_valid_a(array_14_io_d_in_21_valid_a),
    .io_d_in_21_b(array_14_io_d_in_21_b),
    .io_d_in_22_a(array_14_io_d_in_22_a),
    .io_d_in_22_valid_a(array_14_io_d_in_22_valid_a),
    .io_d_in_22_b(array_14_io_d_in_22_b),
    .io_d_in_23_a(array_14_io_d_in_23_a),
    .io_d_in_23_valid_a(array_14_io_d_in_23_valid_a),
    .io_d_in_23_b(array_14_io_d_in_23_b),
    .io_d_in_24_a(array_14_io_d_in_24_a),
    .io_d_in_24_valid_a(array_14_io_d_in_24_valid_a),
    .io_d_in_24_b(array_14_io_d_in_24_b),
    .io_d_in_25_a(array_14_io_d_in_25_a),
    .io_d_in_25_valid_a(array_14_io_d_in_25_valid_a),
    .io_d_in_25_b(array_14_io_d_in_25_b),
    .io_d_in_26_a(array_14_io_d_in_26_a),
    .io_d_in_26_valid_a(array_14_io_d_in_26_valid_a),
    .io_d_in_26_b(array_14_io_d_in_26_b),
    .io_d_in_27_a(array_14_io_d_in_27_a),
    .io_d_in_27_valid_a(array_14_io_d_in_27_valid_a),
    .io_d_in_27_b(array_14_io_d_in_27_b),
    .io_d_in_28_a(array_14_io_d_in_28_a),
    .io_d_in_28_valid_a(array_14_io_d_in_28_valid_a),
    .io_d_in_28_b(array_14_io_d_in_28_b),
    .io_d_in_29_a(array_14_io_d_in_29_a),
    .io_d_in_29_valid_a(array_14_io_d_in_29_valid_a),
    .io_d_in_29_b(array_14_io_d_in_29_b),
    .io_d_in_30_a(array_14_io_d_in_30_a),
    .io_d_in_30_valid_a(array_14_io_d_in_30_valid_a),
    .io_d_in_30_b(array_14_io_d_in_30_b),
    .io_d_in_31_a(array_14_io_d_in_31_a),
    .io_d_in_31_valid_a(array_14_io_d_in_31_valid_a),
    .io_d_in_31_b(array_14_io_d_in_31_b),
    .io_d_out_0_a(array_14_io_d_out_0_a),
    .io_d_out_0_valid_a(array_14_io_d_out_0_valid_a),
    .io_d_out_0_b(array_14_io_d_out_0_b),
    .io_d_out_0_valid_b(array_14_io_d_out_0_valid_b),
    .io_d_out_1_a(array_14_io_d_out_1_a),
    .io_d_out_1_valid_a(array_14_io_d_out_1_valid_a),
    .io_d_out_1_b(array_14_io_d_out_1_b),
    .io_d_out_1_valid_b(array_14_io_d_out_1_valid_b),
    .io_d_out_2_a(array_14_io_d_out_2_a),
    .io_d_out_2_valid_a(array_14_io_d_out_2_valid_a),
    .io_d_out_2_b(array_14_io_d_out_2_b),
    .io_d_out_2_valid_b(array_14_io_d_out_2_valid_b),
    .io_d_out_3_a(array_14_io_d_out_3_a),
    .io_d_out_3_valid_a(array_14_io_d_out_3_valid_a),
    .io_d_out_3_b(array_14_io_d_out_3_b),
    .io_d_out_3_valid_b(array_14_io_d_out_3_valid_b),
    .io_d_out_4_a(array_14_io_d_out_4_a),
    .io_d_out_4_valid_a(array_14_io_d_out_4_valid_a),
    .io_d_out_4_b(array_14_io_d_out_4_b),
    .io_d_out_4_valid_b(array_14_io_d_out_4_valid_b),
    .io_d_out_5_a(array_14_io_d_out_5_a),
    .io_d_out_5_valid_a(array_14_io_d_out_5_valid_a),
    .io_d_out_5_b(array_14_io_d_out_5_b),
    .io_d_out_5_valid_b(array_14_io_d_out_5_valid_b),
    .io_d_out_6_a(array_14_io_d_out_6_a),
    .io_d_out_6_valid_a(array_14_io_d_out_6_valid_a),
    .io_d_out_6_b(array_14_io_d_out_6_b),
    .io_d_out_6_valid_b(array_14_io_d_out_6_valid_b),
    .io_d_out_7_a(array_14_io_d_out_7_a),
    .io_d_out_7_valid_a(array_14_io_d_out_7_valid_a),
    .io_d_out_7_b(array_14_io_d_out_7_b),
    .io_d_out_7_valid_b(array_14_io_d_out_7_valid_b),
    .io_d_out_8_a(array_14_io_d_out_8_a),
    .io_d_out_8_valid_a(array_14_io_d_out_8_valid_a),
    .io_d_out_8_b(array_14_io_d_out_8_b),
    .io_d_out_8_valid_b(array_14_io_d_out_8_valid_b),
    .io_d_out_9_a(array_14_io_d_out_9_a),
    .io_d_out_9_valid_a(array_14_io_d_out_9_valid_a),
    .io_d_out_9_b(array_14_io_d_out_9_b),
    .io_d_out_9_valid_b(array_14_io_d_out_9_valid_b),
    .io_d_out_10_a(array_14_io_d_out_10_a),
    .io_d_out_10_valid_a(array_14_io_d_out_10_valid_a),
    .io_d_out_10_b(array_14_io_d_out_10_b),
    .io_d_out_10_valid_b(array_14_io_d_out_10_valid_b),
    .io_d_out_11_a(array_14_io_d_out_11_a),
    .io_d_out_11_valid_a(array_14_io_d_out_11_valid_a),
    .io_d_out_11_b(array_14_io_d_out_11_b),
    .io_d_out_11_valid_b(array_14_io_d_out_11_valid_b),
    .io_d_out_12_a(array_14_io_d_out_12_a),
    .io_d_out_12_valid_a(array_14_io_d_out_12_valid_a),
    .io_d_out_12_b(array_14_io_d_out_12_b),
    .io_d_out_12_valid_b(array_14_io_d_out_12_valid_b),
    .io_d_out_13_a(array_14_io_d_out_13_a),
    .io_d_out_13_valid_a(array_14_io_d_out_13_valid_a),
    .io_d_out_13_b(array_14_io_d_out_13_b),
    .io_d_out_13_valid_b(array_14_io_d_out_13_valid_b),
    .io_d_out_14_a(array_14_io_d_out_14_a),
    .io_d_out_14_valid_a(array_14_io_d_out_14_valid_a),
    .io_d_out_14_b(array_14_io_d_out_14_b),
    .io_d_out_14_valid_b(array_14_io_d_out_14_valid_b),
    .io_d_out_15_a(array_14_io_d_out_15_a),
    .io_d_out_15_valid_a(array_14_io_d_out_15_valid_a),
    .io_d_out_15_b(array_14_io_d_out_15_b),
    .io_d_out_15_valid_b(array_14_io_d_out_15_valid_b),
    .io_d_out_16_a(array_14_io_d_out_16_a),
    .io_d_out_16_valid_a(array_14_io_d_out_16_valid_a),
    .io_d_out_16_b(array_14_io_d_out_16_b),
    .io_d_out_16_valid_b(array_14_io_d_out_16_valid_b),
    .io_d_out_17_a(array_14_io_d_out_17_a),
    .io_d_out_17_valid_a(array_14_io_d_out_17_valid_a),
    .io_d_out_17_b(array_14_io_d_out_17_b),
    .io_d_out_17_valid_b(array_14_io_d_out_17_valid_b),
    .io_d_out_18_a(array_14_io_d_out_18_a),
    .io_d_out_18_valid_a(array_14_io_d_out_18_valid_a),
    .io_d_out_18_b(array_14_io_d_out_18_b),
    .io_d_out_18_valid_b(array_14_io_d_out_18_valid_b),
    .io_d_out_19_a(array_14_io_d_out_19_a),
    .io_d_out_19_valid_a(array_14_io_d_out_19_valid_a),
    .io_d_out_19_b(array_14_io_d_out_19_b),
    .io_d_out_19_valid_b(array_14_io_d_out_19_valid_b),
    .io_d_out_20_a(array_14_io_d_out_20_a),
    .io_d_out_20_valid_a(array_14_io_d_out_20_valid_a),
    .io_d_out_20_b(array_14_io_d_out_20_b),
    .io_d_out_20_valid_b(array_14_io_d_out_20_valid_b),
    .io_d_out_21_a(array_14_io_d_out_21_a),
    .io_d_out_21_valid_a(array_14_io_d_out_21_valid_a),
    .io_d_out_21_b(array_14_io_d_out_21_b),
    .io_d_out_21_valid_b(array_14_io_d_out_21_valid_b),
    .io_d_out_22_a(array_14_io_d_out_22_a),
    .io_d_out_22_valid_a(array_14_io_d_out_22_valid_a),
    .io_d_out_22_b(array_14_io_d_out_22_b),
    .io_d_out_22_valid_b(array_14_io_d_out_22_valid_b),
    .io_d_out_23_a(array_14_io_d_out_23_a),
    .io_d_out_23_valid_a(array_14_io_d_out_23_valid_a),
    .io_d_out_23_b(array_14_io_d_out_23_b),
    .io_d_out_23_valid_b(array_14_io_d_out_23_valid_b),
    .io_d_out_24_a(array_14_io_d_out_24_a),
    .io_d_out_24_valid_a(array_14_io_d_out_24_valid_a),
    .io_d_out_24_b(array_14_io_d_out_24_b),
    .io_d_out_24_valid_b(array_14_io_d_out_24_valid_b),
    .io_d_out_25_a(array_14_io_d_out_25_a),
    .io_d_out_25_valid_a(array_14_io_d_out_25_valid_a),
    .io_d_out_25_b(array_14_io_d_out_25_b),
    .io_d_out_25_valid_b(array_14_io_d_out_25_valid_b),
    .io_d_out_26_a(array_14_io_d_out_26_a),
    .io_d_out_26_valid_a(array_14_io_d_out_26_valid_a),
    .io_d_out_26_b(array_14_io_d_out_26_b),
    .io_d_out_26_valid_b(array_14_io_d_out_26_valid_b),
    .io_d_out_27_a(array_14_io_d_out_27_a),
    .io_d_out_27_valid_a(array_14_io_d_out_27_valid_a),
    .io_d_out_27_b(array_14_io_d_out_27_b),
    .io_d_out_27_valid_b(array_14_io_d_out_27_valid_b),
    .io_d_out_28_a(array_14_io_d_out_28_a),
    .io_d_out_28_valid_a(array_14_io_d_out_28_valid_a),
    .io_d_out_28_b(array_14_io_d_out_28_b),
    .io_d_out_28_valid_b(array_14_io_d_out_28_valid_b),
    .io_d_out_29_a(array_14_io_d_out_29_a),
    .io_d_out_29_valid_a(array_14_io_d_out_29_valid_a),
    .io_d_out_29_b(array_14_io_d_out_29_b),
    .io_d_out_29_valid_b(array_14_io_d_out_29_valid_b),
    .io_d_out_30_a(array_14_io_d_out_30_a),
    .io_d_out_30_valid_a(array_14_io_d_out_30_valid_a),
    .io_d_out_30_b(array_14_io_d_out_30_b),
    .io_d_out_30_valid_b(array_14_io_d_out_30_valid_b),
    .io_d_out_31_a(array_14_io_d_out_31_a),
    .io_d_out_31_valid_a(array_14_io_d_out_31_valid_a),
    .io_d_out_31_b(array_14_io_d_out_31_b),
    .io_d_out_31_valid_b(array_14_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_14_io_wr_en_mem1),
    .io_wr_en_mem2(array_14_io_wr_en_mem2),
    .io_wr_en_mem3(array_14_io_wr_en_mem3),
    .io_wr_en_mem4(array_14_io_wr_en_mem4),
    .io_wr_en_mem5(array_14_io_wr_en_mem5),
    .io_wr_en_mem6(array_14_io_wr_en_mem6),
    .io_wr_instr_mem1(array_14_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_14_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_14_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_14_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_14_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_14_io_wr_instr_mem6),
    .io_PC1_in(array_14_io_PC1_in),
    .io_PC6_out(array_14_io_PC6_out),
    .io_Addr_in(array_14_io_Addr_in),
    .io_Addr_out(array_14_io_Addr_out),
    .io_Tag_in_Tag(array_14_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_14_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_14_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_14_io_Tag_out_RoundCnt)
  );
  BuildingBlockNew array_15 ( // @[Array.scala 41:54]
    .clock(array_15_clock),
    .reset(array_15_reset),
    .io_d_in_0_a(array_15_io_d_in_0_a),
    .io_d_in_0_valid_a(array_15_io_d_in_0_valid_a),
    .io_d_in_0_b(array_15_io_d_in_0_b),
    .io_d_in_1_a(array_15_io_d_in_1_a),
    .io_d_in_1_valid_a(array_15_io_d_in_1_valid_a),
    .io_d_in_1_b(array_15_io_d_in_1_b),
    .io_d_in_2_a(array_15_io_d_in_2_a),
    .io_d_in_2_valid_a(array_15_io_d_in_2_valid_a),
    .io_d_in_2_b(array_15_io_d_in_2_b),
    .io_d_in_3_a(array_15_io_d_in_3_a),
    .io_d_in_3_valid_a(array_15_io_d_in_3_valid_a),
    .io_d_in_3_b(array_15_io_d_in_3_b),
    .io_d_in_4_a(array_15_io_d_in_4_a),
    .io_d_in_4_valid_a(array_15_io_d_in_4_valid_a),
    .io_d_in_4_b(array_15_io_d_in_4_b),
    .io_d_in_5_a(array_15_io_d_in_5_a),
    .io_d_in_5_valid_a(array_15_io_d_in_5_valid_a),
    .io_d_in_5_b(array_15_io_d_in_5_b),
    .io_d_in_6_a(array_15_io_d_in_6_a),
    .io_d_in_6_valid_a(array_15_io_d_in_6_valid_a),
    .io_d_in_6_b(array_15_io_d_in_6_b),
    .io_d_in_7_a(array_15_io_d_in_7_a),
    .io_d_in_7_valid_a(array_15_io_d_in_7_valid_a),
    .io_d_in_7_b(array_15_io_d_in_7_b),
    .io_d_in_8_a(array_15_io_d_in_8_a),
    .io_d_in_8_valid_a(array_15_io_d_in_8_valid_a),
    .io_d_in_8_b(array_15_io_d_in_8_b),
    .io_d_in_9_a(array_15_io_d_in_9_a),
    .io_d_in_9_valid_a(array_15_io_d_in_9_valid_a),
    .io_d_in_9_b(array_15_io_d_in_9_b),
    .io_d_in_10_a(array_15_io_d_in_10_a),
    .io_d_in_10_valid_a(array_15_io_d_in_10_valid_a),
    .io_d_in_10_b(array_15_io_d_in_10_b),
    .io_d_in_11_a(array_15_io_d_in_11_a),
    .io_d_in_11_valid_a(array_15_io_d_in_11_valid_a),
    .io_d_in_11_b(array_15_io_d_in_11_b),
    .io_d_in_12_a(array_15_io_d_in_12_a),
    .io_d_in_12_valid_a(array_15_io_d_in_12_valid_a),
    .io_d_in_12_b(array_15_io_d_in_12_b),
    .io_d_in_13_a(array_15_io_d_in_13_a),
    .io_d_in_13_valid_a(array_15_io_d_in_13_valid_a),
    .io_d_in_13_b(array_15_io_d_in_13_b),
    .io_d_in_14_a(array_15_io_d_in_14_a),
    .io_d_in_14_valid_a(array_15_io_d_in_14_valid_a),
    .io_d_in_14_b(array_15_io_d_in_14_b),
    .io_d_in_15_a(array_15_io_d_in_15_a),
    .io_d_in_15_valid_a(array_15_io_d_in_15_valid_a),
    .io_d_in_15_b(array_15_io_d_in_15_b),
    .io_d_in_16_a(array_15_io_d_in_16_a),
    .io_d_in_16_valid_a(array_15_io_d_in_16_valid_a),
    .io_d_in_16_b(array_15_io_d_in_16_b),
    .io_d_in_17_a(array_15_io_d_in_17_a),
    .io_d_in_17_valid_a(array_15_io_d_in_17_valid_a),
    .io_d_in_17_b(array_15_io_d_in_17_b),
    .io_d_in_18_a(array_15_io_d_in_18_a),
    .io_d_in_18_valid_a(array_15_io_d_in_18_valid_a),
    .io_d_in_18_b(array_15_io_d_in_18_b),
    .io_d_in_19_a(array_15_io_d_in_19_a),
    .io_d_in_19_valid_a(array_15_io_d_in_19_valid_a),
    .io_d_in_19_b(array_15_io_d_in_19_b),
    .io_d_in_20_a(array_15_io_d_in_20_a),
    .io_d_in_20_valid_a(array_15_io_d_in_20_valid_a),
    .io_d_in_20_b(array_15_io_d_in_20_b),
    .io_d_in_21_a(array_15_io_d_in_21_a),
    .io_d_in_21_valid_a(array_15_io_d_in_21_valid_a),
    .io_d_in_21_b(array_15_io_d_in_21_b),
    .io_d_in_22_a(array_15_io_d_in_22_a),
    .io_d_in_22_valid_a(array_15_io_d_in_22_valid_a),
    .io_d_in_22_b(array_15_io_d_in_22_b),
    .io_d_in_23_a(array_15_io_d_in_23_a),
    .io_d_in_23_valid_a(array_15_io_d_in_23_valid_a),
    .io_d_in_23_b(array_15_io_d_in_23_b),
    .io_d_in_24_a(array_15_io_d_in_24_a),
    .io_d_in_24_valid_a(array_15_io_d_in_24_valid_a),
    .io_d_in_24_b(array_15_io_d_in_24_b),
    .io_d_in_25_a(array_15_io_d_in_25_a),
    .io_d_in_25_valid_a(array_15_io_d_in_25_valid_a),
    .io_d_in_25_b(array_15_io_d_in_25_b),
    .io_d_in_26_a(array_15_io_d_in_26_a),
    .io_d_in_26_valid_a(array_15_io_d_in_26_valid_a),
    .io_d_in_26_b(array_15_io_d_in_26_b),
    .io_d_in_27_a(array_15_io_d_in_27_a),
    .io_d_in_27_valid_a(array_15_io_d_in_27_valid_a),
    .io_d_in_27_b(array_15_io_d_in_27_b),
    .io_d_in_28_a(array_15_io_d_in_28_a),
    .io_d_in_28_valid_a(array_15_io_d_in_28_valid_a),
    .io_d_in_28_b(array_15_io_d_in_28_b),
    .io_d_in_29_a(array_15_io_d_in_29_a),
    .io_d_in_29_valid_a(array_15_io_d_in_29_valid_a),
    .io_d_in_29_b(array_15_io_d_in_29_b),
    .io_d_in_30_a(array_15_io_d_in_30_a),
    .io_d_in_30_valid_a(array_15_io_d_in_30_valid_a),
    .io_d_in_30_b(array_15_io_d_in_30_b),
    .io_d_in_31_a(array_15_io_d_in_31_a),
    .io_d_in_31_valid_a(array_15_io_d_in_31_valid_a),
    .io_d_in_31_b(array_15_io_d_in_31_b),
    .io_d_out_0_a(array_15_io_d_out_0_a),
    .io_d_out_0_valid_a(array_15_io_d_out_0_valid_a),
    .io_d_out_0_b(array_15_io_d_out_0_b),
    .io_d_out_0_valid_b(array_15_io_d_out_0_valid_b),
    .io_d_out_1_a(array_15_io_d_out_1_a),
    .io_d_out_1_valid_a(array_15_io_d_out_1_valid_a),
    .io_d_out_1_b(array_15_io_d_out_1_b),
    .io_d_out_1_valid_b(array_15_io_d_out_1_valid_b),
    .io_d_out_2_a(array_15_io_d_out_2_a),
    .io_d_out_2_valid_a(array_15_io_d_out_2_valid_a),
    .io_d_out_2_b(array_15_io_d_out_2_b),
    .io_d_out_2_valid_b(array_15_io_d_out_2_valid_b),
    .io_d_out_3_a(array_15_io_d_out_3_a),
    .io_d_out_3_valid_a(array_15_io_d_out_3_valid_a),
    .io_d_out_3_b(array_15_io_d_out_3_b),
    .io_d_out_3_valid_b(array_15_io_d_out_3_valid_b),
    .io_d_out_4_a(array_15_io_d_out_4_a),
    .io_d_out_4_valid_a(array_15_io_d_out_4_valid_a),
    .io_d_out_4_b(array_15_io_d_out_4_b),
    .io_d_out_4_valid_b(array_15_io_d_out_4_valid_b),
    .io_d_out_5_a(array_15_io_d_out_5_a),
    .io_d_out_5_valid_a(array_15_io_d_out_5_valid_a),
    .io_d_out_5_b(array_15_io_d_out_5_b),
    .io_d_out_5_valid_b(array_15_io_d_out_5_valid_b),
    .io_d_out_6_a(array_15_io_d_out_6_a),
    .io_d_out_6_valid_a(array_15_io_d_out_6_valid_a),
    .io_d_out_6_b(array_15_io_d_out_6_b),
    .io_d_out_6_valid_b(array_15_io_d_out_6_valid_b),
    .io_d_out_7_a(array_15_io_d_out_7_a),
    .io_d_out_7_valid_a(array_15_io_d_out_7_valid_a),
    .io_d_out_7_b(array_15_io_d_out_7_b),
    .io_d_out_7_valid_b(array_15_io_d_out_7_valid_b),
    .io_d_out_8_a(array_15_io_d_out_8_a),
    .io_d_out_8_valid_a(array_15_io_d_out_8_valid_a),
    .io_d_out_8_b(array_15_io_d_out_8_b),
    .io_d_out_8_valid_b(array_15_io_d_out_8_valid_b),
    .io_d_out_9_a(array_15_io_d_out_9_a),
    .io_d_out_9_valid_a(array_15_io_d_out_9_valid_a),
    .io_d_out_9_b(array_15_io_d_out_9_b),
    .io_d_out_9_valid_b(array_15_io_d_out_9_valid_b),
    .io_d_out_10_a(array_15_io_d_out_10_a),
    .io_d_out_10_valid_a(array_15_io_d_out_10_valid_a),
    .io_d_out_10_b(array_15_io_d_out_10_b),
    .io_d_out_10_valid_b(array_15_io_d_out_10_valid_b),
    .io_d_out_11_a(array_15_io_d_out_11_a),
    .io_d_out_11_valid_a(array_15_io_d_out_11_valid_a),
    .io_d_out_11_b(array_15_io_d_out_11_b),
    .io_d_out_11_valid_b(array_15_io_d_out_11_valid_b),
    .io_d_out_12_a(array_15_io_d_out_12_a),
    .io_d_out_12_valid_a(array_15_io_d_out_12_valid_a),
    .io_d_out_12_b(array_15_io_d_out_12_b),
    .io_d_out_12_valid_b(array_15_io_d_out_12_valid_b),
    .io_d_out_13_a(array_15_io_d_out_13_a),
    .io_d_out_13_valid_a(array_15_io_d_out_13_valid_a),
    .io_d_out_13_b(array_15_io_d_out_13_b),
    .io_d_out_13_valid_b(array_15_io_d_out_13_valid_b),
    .io_d_out_14_a(array_15_io_d_out_14_a),
    .io_d_out_14_valid_a(array_15_io_d_out_14_valid_a),
    .io_d_out_14_b(array_15_io_d_out_14_b),
    .io_d_out_14_valid_b(array_15_io_d_out_14_valid_b),
    .io_d_out_15_a(array_15_io_d_out_15_a),
    .io_d_out_15_valid_a(array_15_io_d_out_15_valid_a),
    .io_d_out_15_b(array_15_io_d_out_15_b),
    .io_d_out_15_valid_b(array_15_io_d_out_15_valid_b),
    .io_d_out_16_a(array_15_io_d_out_16_a),
    .io_d_out_16_valid_a(array_15_io_d_out_16_valid_a),
    .io_d_out_16_b(array_15_io_d_out_16_b),
    .io_d_out_16_valid_b(array_15_io_d_out_16_valid_b),
    .io_d_out_17_a(array_15_io_d_out_17_a),
    .io_d_out_17_valid_a(array_15_io_d_out_17_valid_a),
    .io_d_out_17_b(array_15_io_d_out_17_b),
    .io_d_out_17_valid_b(array_15_io_d_out_17_valid_b),
    .io_d_out_18_a(array_15_io_d_out_18_a),
    .io_d_out_18_valid_a(array_15_io_d_out_18_valid_a),
    .io_d_out_18_b(array_15_io_d_out_18_b),
    .io_d_out_18_valid_b(array_15_io_d_out_18_valid_b),
    .io_d_out_19_a(array_15_io_d_out_19_a),
    .io_d_out_19_valid_a(array_15_io_d_out_19_valid_a),
    .io_d_out_19_b(array_15_io_d_out_19_b),
    .io_d_out_19_valid_b(array_15_io_d_out_19_valid_b),
    .io_d_out_20_a(array_15_io_d_out_20_a),
    .io_d_out_20_valid_a(array_15_io_d_out_20_valid_a),
    .io_d_out_20_b(array_15_io_d_out_20_b),
    .io_d_out_20_valid_b(array_15_io_d_out_20_valid_b),
    .io_d_out_21_a(array_15_io_d_out_21_a),
    .io_d_out_21_valid_a(array_15_io_d_out_21_valid_a),
    .io_d_out_21_b(array_15_io_d_out_21_b),
    .io_d_out_21_valid_b(array_15_io_d_out_21_valid_b),
    .io_d_out_22_a(array_15_io_d_out_22_a),
    .io_d_out_22_valid_a(array_15_io_d_out_22_valid_a),
    .io_d_out_22_b(array_15_io_d_out_22_b),
    .io_d_out_22_valid_b(array_15_io_d_out_22_valid_b),
    .io_d_out_23_a(array_15_io_d_out_23_a),
    .io_d_out_23_valid_a(array_15_io_d_out_23_valid_a),
    .io_d_out_23_b(array_15_io_d_out_23_b),
    .io_d_out_23_valid_b(array_15_io_d_out_23_valid_b),
    .io_d_out_24_a(array_15_io_d_out_24_a),
    .io_d_out_24_valid_a(array_15_io_d_out_24_valid_a),
    .io_d_out_24_b(array_15_io_d_out_24_b),
    .io_d_out_24_valid_b(array_15_io_d_out_24_valid_b),
    .io_d_out_25_a(array_15_io_d_out_25_a),
    .io_d_out_25_valid_a(array_15_io_d_out_25_valid_a),
    .io_d_out_25_b(array_15_io_d_out_25_b),
    .io_d_out_25_valid_b(array_15_io_d_out_25_valid_b),
    .io_d_out_26_a(array_15_io_d_out_26_a),
    .io_d_out_26_valid_a(array_15_io_d_out_26_valid_a),
    .io_d_out_26_b(array_15_io_d_out_26_b),
    .io_d_out_26_valid_b(array_15_io_d_out_26_valid_b),
    .io_d_out_27_a(array_15_io_d_out_27_a),
    .io_d_out_27_valid_a(array_15_io_d_out_27_valid_a),
    .io_d_out_27_b(array_15_io_d_out_27_b),
    .io_d_out_27_valid_b(array_15_io_d_out_27_valid_b),
    .io_d_out_28_a(array_15_io_d_out_28_a),
    .io_d_out_28_valid_a(array_15_io_d_out_28_valid_a),
    .io_d_out_28_b(array_15_io_d_out_28_b),
    .io_d_out_28_valid_b(array_15_io_d_out_28_valid_b),
    .io_d_out_29_a(array_15_io_d_out_29_a),
    .io_d_out_29_valid_a(array_15_io_d_out_29_valid_a),
    .io_d_out_29_b(array_15_io_d_out_29_b),
    .io_d_out_29_valid_b(array_15_io_d_out_29_valid_b),
    .io_d_out_30_a(array_15_io_d_out_30_a),
    .io_d_out_30_valid_a(array_15_io_d_out_30_valid_a),
    .io_d_out_30_b(array_15_io_d_out_30_b),
    .io_d_out_30_valid_b(array_15_io_d_out_30_valid_b),
    .io_d_out_31_a(array_15_io_d_out_31_a),
    .io_d_out_31_valid_a(array_15_io_d_out_31_valid_a),
    .io_d_out_31_b(array_15_io_d_out_31_b),
    .io_d_out_31_valid_b(array_15_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_15_io_wr_en_mem1),
    .io_wr_en_mem2(array_15_io_wr_en_mem2),
    .io_wr_en_mem3(array_15_io_wr_en_mem3),
    .io_wr_en_mem4(array_15_io_wr_en_mem4),
    .io_wr_en_mem5(array_15_io_wr_en_mem5),
    .io_wr_en_mem6(array_15_io_wr_en_mem6),
    .io_wr_instr_mem1(array_15_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_15_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_15_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_15_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_15_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_15_io_wr_instr_mem6),
    .io_PC1_in(array_15_io_PC1_in),
    .io_PC6_out(array_15_io_PC6_out),
    .io_Addr_in(array_15_io_Addr_in),
    .io_Addr_out(array_15_io_Addr_out),
    .io_Tag_in_Tag(array_15_io_Tag_in_Tag),
    .io_Tag_in_RoundCnt(array_15_io_Tag_in_RoundCnt),
    .io_Tag_out_Tag(array_15_io_Tag_out_Tag),
    .io_Tag_out_RoundCnt(array_15_io_Tag_out_RoundCnt)
  );
  assign io_d_out_0_a = array_15_io_d_out_0_a; // @[Array.scala 88:12]
  assign io_d_out_0_valid_a = array_15_io_d_out_0_valid_a; // @[Array.scala 88:12]
  assign io_d_out_0_b = array_15_io_d_out_0_b; // @[Array.scala 88:12]
  assign io_d_out_0_valid_b = array_15_io_d_out_0_valid_b; // @[Array.scala 88:12]
  assign io_d_out_1_a = array_15_io_d_out_1_a; // @[Array.scala 88:12]
  assign io_d_out_1_valid_a = array_15_io_d_out_1_valid_a; // @[Array.scala 88:12]
  assign io_d_out_1_b = array_15_io_d_out_1_b; // @[Array.scala 88:12]
  assign io_d_out_1_valid_b = array_15_io_d_out_1_valid_b; // @[Array.scala 88:12]
  assign io_d_out_2_a = array_15_io_d_out_2_a; // @[Array.scala 88:12]
  assign io_d_out_2_valid_a = array_15_io_d_out_2_valid_a; // @[Array.scala 88:12]
  assign io_d_out_2_b = array_15_io_d_out_2_b; // @[Array.scala 88:12]
  assign io_d_out_2_valid_b = array_15_io_d_out_2_valid_b; // @[Array.scala 88:12]
  assign io_d_out_3_a = array_15_io_d_out_3_a; // @[Array.scala 88:12]
  assign io_d_out_3_valid_a = array_15_io_d_out_3_valid_a; // @[Array.scala 88:12]
  assign io_d_out_3_b = array_15_io_d_out_3_b; // @[Array.scala 88:12]
  assign io_d_out_3_valid_b = array_15_io_d_out_3_valid_b; // @[Array.scala 88:12]
  assign io_d_out_4_a = array_15_io_d_out_4_a; // @[Array.scala 88:12]
  assign io_d_out_4_valid_a = array_15_io_d_out_4_valid_a; // @[Array.scala 88:12]
  assign io_d_out_4_b = array_15_io_d_out_4_b; // @[Array.scala 88:12]
  assign io_d_out_4_valid_b = array_15_io_d_out_4_valid_b; // @[Array.scala 88:12]
  assign io_d_out_5_a = array_15_io_d_out_5_a; // @[Array.scala 88:12]
  assign io_d_out_5_valid_a = array_15_io_d_out_5_valid_a; // @[Array.scala 88:12]
  assign io_d_out_5_b = array_15_io_d_out_5_b; // @[Array.scala 88:12]
  assign io_d_out_5_valid_b = array_15_io_d_out_5_valid_b; // @[Array.scala 88:12]
  assign io_d_out_6_a = array_15_io_d_out_6_a; // @[Array.scala 88:12]
  assign io_d_out_6_valid_a = array_15_io_d_out_6_valid_a; // @[Array.scala 88:12]
  assign io_d_out_6_b = array_15_io_d_out_6_b; // @[Array.scala 88:12]
  assign io_d_out_6_valid_b = array_15_io_d_out_6_valid_b; // @[Array.scala 88:12]
  assign io_d_out_7_a = array_15_io_d_out_7_a; // @[Array.scala 88:12]
  assign io_d_out_7_valid_a = array_15_io_d_out_7_valid_a; // @[Array.scala 88:12]
  assign io_d_out_7_b = array_15_io_d_out_7_b; // @[Array.scala 88:12]
  assign io_d_out_7_valid_b = array_15_io_d_out_7_valid_b; // @[Array.scala 88:12]
  assign io_d_out_8_a = array_15_io_d_out_8_a; // @[Array.scala 88:12]
  assign io_d_out_8_valid_a = array_15_io_d_out_8_valid_a; // @[Array.scala 88:12]
  assign io_d_out_8_b = array_15_io_d_out_8_b; // @[Array.scala 88:12]
  assign io_d_out_8_valid_b = array_15_io_d_out_8_valid_b; // @[Array.scala 88:12]
  assign io_d_out_9_a = array_15_io_d_out_9_a; // @[Array.scala 88:12]
  assign io_d_out_9_valid_a = array_15_io_d_out_9_valid_a; // @[Array.scala 88:12]
  assign io_d_out_9_b = array_15_io_d_out_9_b; // @[Array.scala 88:12]
  assign io_d_out_9_valid_b = array_15_io_d_out_9_valid_b; // @[Array.scala 88:12]
  assign io_d_out_10_a = array_15_io_d_out_10_a; // @[Array.scala 88:12]
  assign io_d_out_10_valid_a = array_15_io_d_out_10_valid_a; // @[Array.scala 88:12]
  assign io_d_out_10_b = array_15_io_d_out_10_b; // @[Array.scala 88:12]
  assign io_d_out_10_valid_b = array_15_io_d_out_10_valid_b; // @[Array.scala 88:12]
  assign io_d_out_11_a = array_15_io_d_out_11_a; // @[Array.scala 88:12]
  assign io_d_out_11_valid_a = array_15_io_d_out_11_valid_a; // @[Array.scala 88:12]
  assign io_d_out_11_b = array_15_io_d_out_11_b; // @[Array.scala 88:12]
  assign io_d_out_11_valid_b = array_15_io_d_out_11_valid_b; // @[Array.scala 88:12]
  assign io_d_out_12_a = array_15_io_d_out_12_a; // @[Array.scala 88:12]
  assign io_d_out_12_valid_a = array_15_io_d_out_12_valid_a; // @[Array.scala 88:12]
  assign io_d_out_12_b = array_15_io_d_out_12_b; // @[Array.scala 88:12]
  assign io_d_out_12_valid_b = array_15_io_d_out_12_valid_b; // @[Array.scala 88:12]
  assign io_d_out_13_a = array_15_io_d_out_13_a; // @[Array.scala 88:12]
  assign io_d_out_13_valid_a = array_15_io_d_out_13_valid_a; // @[Array.scala 88:12]
  assign io_d_out_13_b = array_15_io_d_out_13_b; // @[Array.scala 88:12]
  assign io_d_out_13_valid_b = array_15_io_d_out_13_valid_b; // @[Array.scala 88:12]
  assign io_d_out_14_a = array_15_io_d_out_14_a; // @[Array.scala 88:12]
  assign io_d_out_14_valid_a = array_15_io_d_out_14_valid_a; // @[Array.scala 88:12]
  assign io_d_out_14_b = array_15_io_d_out_14_b; // @[Array.scala 88:12]
  assign io_d_out_14_valid_b = array_15_io_d_out_14_valid_b; // @[Array.scala 88:12]
  assign io_d_out_15_a = array_15_io_d_out_15_a; // @[Array.scala 88:12]
  assign io_d_out_15_valid_a = array_15_io_d_out_15_valid_a; // @[Array.scala 88:12]
  assign io_d_out_15_b = array_15_io_d_out_15_b; // @[Array.scala 88:12]
  assign io_d_out_15_valid_b = array_15_io_d_out_15_valid_b; // @[Array.scala 88:12]
  assign io_d_out_16_a = array_15_io_d_out_16_a; // @[Array.scala 88:12]
  assign io_d_out_16_valid_a = array_15_io_d_out_16_valid_a; // @[Array.scala 88:12]
  assign io_d_out_16_b = array_15_io_d_out_16_b; // @[Array.scala 88:12]
  assign io_d_out_16_valid_b = array_15_io_d_out_16_valid_b; // @[Array.scala 88:12]
  assign io_d_out_17_a = array_15_io_d_out_17_a; // @[Array.scala 88:12]
  assign io_d_out_17_valid_a = array_15_io_d_out_17_valid_a; // @[Array.scala 88:12]
  assign io_d_out_17_b = array_15_io_d_out_17_b; // @[Array.scala 88:12]
  assign io_d_out_17_valid_b = array_15_io_d_out_17_valid_b; // @[Array.scala 88:12]
  assign io_d_out_18_a = array_15_io_d_out_18_a; // @[Array.scala 88:12]
  assign io_d_out_18_valid_a = array_15_io_d_out_18_valid_a; // @[Array.scala 88:12]
  assign io_d_out_18_b = array_15_io_d_out_18_b; // @[Array.scala 88:12]
  assign io_d_out_18_valid_b = array_15_io_d_out_18_valid_b; // @[Array.scala 88:12]
  assign io_d_out_19_a = array_15_io_d_out_19_a; // @[Array.scala 88:12]
  assign io_d_out_19_valid_a = array_15_io_d_out_19_valid_a; // @[Array.scala 88:12]
  assign io_d_out_19_b = array_15_io_d_out_19_b; // @[Array.scala 88:12]
  assign io_d_out_19_valid_b = array_15_io_d_out_19_valid_b; // @[Array.scala 88:12]
  assign io_d_out_20_a = array_15_io_d_out_20_a; // @[Array.scala 88:12]
  assign io_d_out_20_valid_a = array_15_io_d_out_20_valid_a; // @[Array.scala 88:12]
  assign io_d_out_20_b = array_15_io_d_out_20_b; // @[Array.scala 88:12]
  assign io_d_out_20_valid_b = array_15_io_d_out_20_valid_b; // @[Array.scala 88:12]
  assign io_d_out_21_a = array_15_io_d_out_21_a; // @[Array.scala 88:12]
  assign io_d_out_21_valid_a = array_15_io_d_out_21_valid_a; // @[Array.scala 88:12]
  assign io_d_out_21_b = array_15_io_d_out_21_b; // @[Array.scala 88:12]
  assign io_d_out_21_valid_b = array_15_io_d_out_21_valid_b; // @[Array.scala 88:12]
  assign io_d_out_22_a = array_15_io_d_out_22_a; // @[Array.scala 88:12]
  assign io_d_out_22_valid_a = array_15_io_d_out_22_valid_a; // @[Array.scala 88:12]
  assign io_d_out_22_b = array_15_io_d_out_22_b; // @[Array.scala 88:12]
  assign io_d_out_22_valid_b = array_15_io_d_out_22_valid_b; // @[Array.scala 88:12]
  assign io_d_out_23_a = array_15_io_d_out_23_a; // @[Array.scala 88:12]
  assign io_d_out_23_valid_a = array_15_io_d_out_23_valid_a; // @[Array.scala 88:12]
  assign io_d_out_23_b = array_15_io_d_out_23_b; // @[Array.scala 88:12]
  assign io_d_out_23_valid_b = array_15_io_d_out_23_valid_b; // @[Array.scala 88:12]
  assign io_d_out_24_a = array_15_io_d_out_24_a; // @[Array.scala 88:12]
  assign io_d_out_24_valid_a = array_15_io_d_out_24_valid_a; // @[Array.scala 88:12]
  assign io_d_out_24_b = array_15_io_d_out_24_b; // @[Array.scala 88:12]
  assign io_d_out_24_valid_b = array_15_io_d_out_24_valid_b; // @[Array.scala 88:12]
  assign io_d_out_25_a = array_15_io_d_out_25_a; // @[Array.scala 88:12]
  assign io_d_out_25_valid_a = array_15_io_d_out_25_valid_a; // @[Array.scala 88:12]
  assign io_d_out_25_b = array_15_io_d_out_25_b; // @[Array.scala 88:12]
  assign io_d_out_25_valid_b = array_15_io_d_out_25_valid_b; // @[Array.scala 88:12]
  assign io_d_out_26_a = array_15_io_d_out_26_a; // @[Array.scala 88:12]
  assign io_d_out_26_valid_a = array_15_io_d_out_26_valid_a; // @[Array.scala 88:12]
  assign io_d_out_26_b = array_15_io_d_out_26_b; // @[Array.scala 88:12]
  assign io_d_out_26_valid_b = array_15_io_d_out_26_valid_b; // @[Array.scala 88:12]
  assign io_d_out_27_a = array_15_io_d_out_27_a; // @[Array.scala 88:12]
  assign io_d_out_27_valid_a = array_15_io_d_out_27_valid_a; // @[Array.scala 88:12]
  assign io_d_out_27_b = array_15_io_d_out_27_b; // @[Array.scala 88:12]
  assign io_d_out_27_valid_b = array_15_io_d_out_27_valid_b; // @[Array.scala 88:12]
  assign io_d_out_28_a = array_15_io_d_out_28_a; // @[Array.scala 88:12]
  assign io_d_out_28_valid_a = array_15_io_d_out_28_valid_a; // @[Array.scala 88:12]
  assign io_d_out_28_b = array_15_io_d_out_28_b; // @[Array.scala 88:12]
  assign io_d_out_28_valid_b = array_15_io_d_out_28_valid_b; // @[Array.scala 88:12]
  assign io_d_out_29_a = array_15_io_d_out_29_a; // @[Array.scala 88:12]
  assign io_d_out_29_valid_a = array_15_io_d_out_29_valid_a; // @[Array.scala 88:12]
  assign io_d_out_29_b = array_15_io_d_out_29_b; // @[Array.scala 88:12]
  assign io_d_out_29_valid_b = array_15_io_d_out_29_valid_b; // @[Array.scala 88:12]
  assign io_d_out_30_a = array_15_io_d_out_30_a; // @[Array.scala 88:12]
  assign io_d_out_30_valid_a = array_15_io_d_out_30_valid_a; // @[Array.scala 88:12]
  assign io_d_out_30_b = array_15_io_d_out_30_b; // @[Array.scala 88:12]
  assign io_d_out_30_valid_b = array_15_io_d_out_30_valid_b; // @[Array.scala 88:12]
  assign io_d_out_31_a = array_15_io_d_out_31_a; // @[Array.scala 88:12]
  assign io_d_out_31_valid_a = array_15_io_d_out_31_valid_a; // @[Array.scala 88:12]
  assign io_d_out_31_b = array_15_io_d_out_31_b; // @[Array.scala 88:12]
  assign io_d_out_31_valid_b = array_15_io_d_out_31_valid_b; // @[Array.scala 88:12]
  assign io_Tag_out_Tag = array_15_io_Tag_out_Tag; // @[Array.scala 89:14]
  assign io_Tag_out_RoundCnt = array_15_io_Tag_out_RoundCnt; // @[Array.scala 89:14]
  assign io_Addr_out = array_15_io_Addr_out; // @[Array.scala 90:15]
  assign io_PC_out = array_15_io_PC6_out; // @[Array.scala 91:13]
  assign array_0_clock = clock;
  assign array_0_reset = reset;
  assign array_0_io_d_in_0_a = io_d_in_0_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_0_valid_a = io_d_in_0_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_0_b = io_d_in_0_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_1_a = io_d_in_1_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_1_valid_a = io_d_in_1_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_1_b = io_d_in_1_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_2_a = io_d_in_2_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_2_valid_a = io_d_in_2_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_2_b = io_d_in_2_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_3_a = io_d_in_3_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_3_valid_a = io_d_in_3_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_3_b = io_d_in_3_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_4_a = io_d_in_4_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_4_valid_a = io_d_in_4_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_4_b = io_d_in_4_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_5_a = io_d_in_5_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_5_valid_a = io_d_in_5_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_5_b = io_d_in_5_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_6_a = io_d_in_6_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_6_valid_a = io_d_in_6_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_6_b = io_d_in_6_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_7_a = io_d_in_7_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_7_valid_a = io_d_in_7_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_7_b = io_d_in_7_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_8_a = io_d_in_8_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_8_valid_a = io_d_in_8_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_8_b = io_d_in_8_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_9_a = io_d_in_9_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_9_valid_a = io_d_in_9_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_9_b = io_d_in_9_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_10_a = io_d_in_10_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_10_valid_a = io_d_in_10_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_10_b = io_d_in_10_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_11_a = io_d_in_11_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_11_valid_a = io_d_in_11_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_11_b = io_d_in_11_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_12_a = io_d_in_12_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_12_valid_a = io_d_in_12_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_12_b = io_d_in_12_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_13_a = io_d_in_13_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_13_valid_a = io_d_in_13_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_13_b = io_d_in_13_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_14_a = io_d_in_14_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_14_valid_a = io_d_in_14_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_14_b = io_d_in_14_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_15_a = io_d_in_15_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_15_valid_a = io_d_in_15_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_15_b = io_d_in_15_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_16_a = io_d_in_16_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_16_valid_a = io_d_in_16_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_16_b = io_d_in_16_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_17_a = io_d_in_17_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_17_valid_a = io_d_in_17_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_17_b = io_d_in_17_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_18_a = io_d_in_18_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_18_valid_a = io_d_in_18_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_18_b = io_d_in_18_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_19_a = io_d_in_19_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_19_valid_a = io_d_in_19_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_19_b = io_d_in_19_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_20_a = io_d_in_20_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_20_valid_a = io_d_in_20_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_20_b = io_d_in_20_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_21_a = io_d_in_21_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_21_valid_a = io_d_in_21_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_21_b = io_d_in_21_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_22_a = io_d_in_22_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_22_valid_a = io_d_in_22_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_22_b = io_d_in_22_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_23_a = io_d_in_23_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_23_valid_a = io_d_in_23_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_23_b = io_d_in_23_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_24_a = io_d_in_24_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_24_valid_a = io_d_in_24_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_24_b = io_d_in_24_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_25_a = io_d_in_25_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_25_valid_a = io_d_in_25_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_25_b = io_d_in_25_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_26_a = io_d_in_26_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_26_valid_a = io_d_in_26_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_26_b = io_d_in_26_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_27_a = io_d_in_27_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_27_valid_a = io_d_in_27_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_27_b = io_d_in_27_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_28_a = io_d_in_28_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_28_valid_a = io_d_in_28_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_28_b = io_d_in_28_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_29_a = io_d_in_29_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_29_valid_a = io_d_in_29_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_29_b = io_d_in_29_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_30_a = io_d_in_30_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_30_valid_a = io_d_in_30_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_30_b = io_d_in_30_b; // @[Array.scala 42:20]
  assign array_0_io_d_in_31_a = io_d_in_31_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_31_valid_a = io_d_in_31_valid_a; // @[Array.scala 42:20]
  assign array_0_io_d_in_31_b = io_d_in_31_b; // @[Array.scala 42:20]
  assign array_0_io_wr_en_mem1 = io_wr_en_mem1_0; // @[Array.scala 52:26]
  assign array_0_io_wr_en_mem2 = io_wr_en_mem2_0; // @[Array.scala 53:26]
  assign array_0_io_wr_en_mem3 = io_wr_en_mem3_0; // @[Array.scala 54:26]
  assign array_0_io_wr_en_mem4 = io_wr_en_mem4_0; // @[Array.scala 55:26]
  assign array_0_io_wr_en_mem5 = io_wr_en_mem5_0; // @[Array.scala 56:26]
  assign array_0_io_wr_en_mem6 = io_wr_en_mem6_0; // @[Array.scala 57:26]
  assign array_0_io_wr_instr_mem1 = io_wr_instr_mem1_0; // @[Array.scala 58:29]
  assign array_0_io_wr_instr_mem2 = io_wr_instr_mem2_0; // @[Array.scala 59:29]
  assign array_0_io_wr_instr_mem3 = io_wr_instr_mem3_0; // @[Array.scala 60:29]
  assign array_0_io_wr_instr_mem4 = io_wr_instr_mem4_0; // @[Array.scala 61:29]
  assign array_0_io_wr_instr_mem5 = io_wr_instr_mem5_0; // @[Array.scala 62:29]
  assign array_0_io_wr_instr_mem6 = io_wr_instr_mem6_0; // @[Array.scala 63:29]
  assign array_0_io_PC1_in = io_PC_in; // @[Array.scala 47:22]
  assign array_0_io_Addr_in = io_Addr_in; // @[Array.scala 48:23]
  assign array_0_io_Tag_in_Tag = io_Tag_in_Tag; // @[Array.scala 43:22]
  assign array_0_io_Tag_in_RoundCnt = io_Tag_in_RoundCnt; // @[Array.scala 43:22]
  assign array_1_clock = clock;
  assign array_1_reset = reset;
  assign array_1_io_d_in_0_a = array_0_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_0_valid_a = array_0_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_0_b = array_0_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_1_a = array_0_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_1_valid_a = array_0_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_1_b = array_0_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_2_a = array_0_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_2_valid_a = array_0_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_2_b = array_0_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_3_a = array_0_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_3_valid_a = array_0_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_3_b = array_0_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_4_a = array_0_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_4_valid_a = array_0_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_4_b = array_0_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_5_a = array_0_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_5_valid_a = array_0_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_5_b = array_0_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_6_a = array_0_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_6_valid_a = array_0_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_6_b = array_0_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_7_a = array_0_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_7_valid_a = array_0_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_7_b = array_0_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_8_a = array_0_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_8_valid_a = array_0_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_8_b = array_0_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_9_a = array_0_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_9_valid_a = array_0_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_9_b = array_0_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_10_a = array_0_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_10_valid_a = array_0_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_10_b = array_0_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_11_a = array_0_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_11_valid_a = array_0_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_11_b = array_0_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_12_a = array_0_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_12_valid_a = array_0_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_12_b = array_0_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_13_a = array_0_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_13_valid_a = array_0_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_13_b = array_0_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_14_a = array_0_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_14_valid_a = array_0_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_14_b = array_0_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_15_a = array_0_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_15_valid_a = array_0_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_15_b = array_0_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_16_a = array_0_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_16_valid_a = array_0_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_16_b = array_0_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_17_a = array_0_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_17_valid_a = array_0_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_17_b = array_0_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_18_a = array_0_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_18_valid_a = array_0_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_18_b = array_0_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_19_a = array_0_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_19_valid_a = array_0_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_19_b = array_0_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_20_a = array_0_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_20_valid_a = array_0_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_20_b = array_0_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_21_a = array_0_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_21_valid_a = array_0_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_21_b = array_0_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_22_a = array_0_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_22_valid_a = array_0_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_22_b = array_0_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_23_a = array_0_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_23_valid_a = array_0_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_23_b = array_0_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_24_a = array_0_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_24_valid_a = array_0_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_24_b = array_0_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_25_a = array_0_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_25_valid_a = array_0_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_25_b = array_0_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_26_a = array_0_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_26_valid_a = array_0_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_26_b = array_0_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_27_a = array_0_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_27_valid_a = array_0_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_27_b = array_0_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_28_a = array_0_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_28_valid_a = array_0_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_28_b = array_0_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_29_a = array_0_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_29_valid_a = array_0_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_29_b = array_0_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_30_a = array_0_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_30_valid_a = array_0_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_30_b = array_0_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_1_io_d_in_31_a = array_0_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_31_valid_a = array_0_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_1_io_d_in_31_b = array_0_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_1_io_wr_en_mem1 = io_wr_en_mem1_1; // @[Array.scala 71:28]
  assign array_1_io_wr_en_mem2 = io_wr_en_mem2_1; // @[Array.scala 72:28]
  assign array_1_io_wr_en_mem3 = io_wr_en_mem3_1; // @[Array.scala 73:28]
  assign array_1_io_wr_en_mem4 = io_wr_en_mem4_1; // @[Array.scala 74:28]
  assign array_1_io_wr_en_mem5 = io_wr_en_mem5_1; // @[Array.scala 75:28]
  assign array_1_io_wr_en_mem6 = io_wr_en_mem6_1; // @[Array.scala 76:28]
  assign array_1_io_wr_instr_mem1 = io_wr_instr_mem1_1; // @[Array.scala 77:31]
  assign array_1_io_wr_instr_mem2 = io_wr_instr_mem2_1; // @[Array.scala 78:31]
  assign array_1_io_wr_instr_mem3 = io_wr_instr_mem3_1; // @[Array.scala 79:31]
  assign array_1_io_wr_instr_mem4 = io_wr_instr_mem4_1; // @[Array.scala 80:31]
  assign array_1_io_wr_instr_mem5 = io_wr_instr_mem5_1; // @[Array.scala 81:31]
  assign array_1_io_wr_instr_mem6 = io_wr_instr_mem6_1; // @[Array.scala 82:31]
  assign array_1_io_PC1_in = array_0_io_PC6_out; // @[Array.scala 84:24]
  assign array_1_io_Addr_in = array_0_io_Addr_out; // @[Array.scala 85:25]
  assign array_1_io_Tag_in_Tag = array_0_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_1_io_Tag_in_RoundCnt = array_0_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
  assign array_2_clock = clock;
  assign array_2_reset = reset;
  assign array_2_io_d_in_0_a = array_1_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_0_valid_a = array_1_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_0_b = array_1_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_1_a = array_1_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_1_valid_a = array_1_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_1_b = array_1_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_2_a = array_1_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_2_valid_a = array_1_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_2_b = array_1_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_3_a = array_1_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_3_valid_a = array_1_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_3_b = array_1_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_4_a = array_1_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_4_valid_a = array_1_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_4_b = array_1_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_5_a = array_1_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_5_valid_a = array_1_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_5_b = array_1_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_6_a = array_1_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_6_valid_a = array_1_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_6_b = array_1_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_7_a = array_1_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_7_valid_a = array_1_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_7_b = array_1_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_8_a = array_1_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_8_valid_a = array_1_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_8_b = array_1_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_9_a = array_1_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_9_valid_a = array_1_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_9_b = array_1_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_10_a = array_1_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_10_valid_a = array_1_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_10_b = array_1_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_11_a = array_1_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_11_valid_a = array_1_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_11_b = array_1_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_12_a = array_1_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_12_valid_a = array_1_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_12_b = array_1_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_13_a = array_1_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_13_valid_a = array_1_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_13_b = array_1_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_14_a = array_1_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_14_valid_a = array_1_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_14_b = array_1_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_15_a = array_1_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_15_valid_a = array_1_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_15_b = array_1_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_16_a = array_1_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_16_valid_a = array_1_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_16_b = array_1_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_17_a = array_1_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_17_valid_a = array_1_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_17_b = array_1_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_18_a = array_1_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_18_valid_a = array_1_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_18_b = array_1_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_19_a = array_1_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_19_valid_a = array_1_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_19_b = array_1_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_20_a = array_1_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_20_valid_a = array_1_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_20_b = array_1_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_21_a = array_1_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_21_valid_a = array_1_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_21_b = array_1_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_22_a = array_1_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_22_valid_a = array_1_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_22_b = array_1_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_23_a = array_1_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_23_valid_a = array_1_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_23_b = array_1_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_24_a = array_1_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_24_valid_a = array_1_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_24_b = array_1_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_25_a = array_1_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_25_valid_a = array_1_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_25_b = array_1_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_26_a = array_1_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_26_valid_a = array_1_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_26_b = array_1_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_27_a = array_1_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_27_valid_a = array_1_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_27_b = array_1_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_28_a = array_1_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_28_valid_a = array_1_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_28_b = array_1_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_29_a = array_1_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_29_valid_a = array_1_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_29_b = array_1_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_30_a = array_1_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_30_valid_a = array_1_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_30_b = array_1_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_2_io_d_in_31_a = array_1_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_31_valid_a = array_1_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_2_io_d_in_31_b = array_1_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_2_io_wr_en_mem1 = io_wr_en_mem1_2; // @[Array.scala 71:28]
  assign array_2_io_wr_en_mem2 = io_wr_en_mem2_2; // @[Array.scala 72:28]
  assign array_2_io_wr_en_mem3 = io_wr_en_mem3_2; // @[Array.scala 73:28]
  assign array_2_io_wr_en_mem4 = io_wr_en_mem4_2; // @[Array.scala 74:28]
  assign array_2_io_wr_en_mem5 = io_wr_en_mem5_2; // @[Array.scala 75:28]
  assign array_2_io_wr_en_mem6 = io_wr_en_mem6_2; // @[Array.scala 76:28]
  assign array_2_io_wr_instr_mem1 = io_wr_instr_mem1_2; // @[Array.scala 77:31]
  assign array_2_io_wr_instr_mem2 = io_wr_instr_mem2_2; // @[Array.scala 78:31]
  assign array_2_io_wr_instr_mem3 = io_wr_instr_mem3_2; // @[Array.scala 79:31]
  assign array_2_io_wr_instr_mem4 = io_wr_instr_mem4_2; // @[Array.scala 80:31]
  assign array_2_io_wr_instr_mem5 = io_wr_instr_mem5_2; // @[Array.scala 81:31]
  assign array_2_io_wr_instr_mem6 = io_wr_instr_mem6_2; // @[Array.scala 82:31]
  assign array_2_io_PC1_in = array_1_io_PC6_out; // @[Array.scala 84:24]
  assign array_2_io_Addr_in = array_1_io_Addr_out; // @[Array.scala 85:25]
  assign array_2_io_Tag_in_Tag = array_1_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_2_io_Tag_in_RoundCnt = array_1_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
  assign array_3_clock = clock;
  assign array_3_reset = reset;
  assign array_3_io_d_in_0_a = array_2_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_0_valid_a = array_2_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_0_b = array_2_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_1_a = array_2_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_1_valid_a = array_2_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_1_b = array_2_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_2_a = array_2_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_2_valid_a = array_2_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_2_b = array_2_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_3_a = array_2_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_3_valid_a = array_2_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_3_b = array_2_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_4_a = array_2_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_4_valid_a = array_2_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_4_b = array_2_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_5_a = array_2_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_5_valid_a = array_2_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_5_b = array_2_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_6_a = array_2_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_6_valid_a = array_2_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_6_b = array_2_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_7_a = array_2_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_7_valid_a = array_2_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_7_b = array_2_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_8_a = array_2_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_8_valid_a = array_2_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_8_b = array_2_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_9_a = array_2_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_9_valid_a = array_2_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_9_b = array_2_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_10_a = array_2_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_10_valid_a = array_2_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_10_b = array_2_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_11_a = array_2_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_11_valid_a = array_2_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_11_b = array_2_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_12_a = array_2_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_12_valid_a = array_2_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_12_b = array_2_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_13_a = array_2_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_13_valid_a = array_2_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_13_b = array_2_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_14_a = array_2_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_14_valid_a = array_2_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_14_b = array_2_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_15_a = array_2_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_15_valid_a = array_2_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_15_b = array_2_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_16_a = array_2_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_16_valid_a = array_2_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_16_b = array_2_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_17_a = array_2_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_17_valid_a = array_2_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_17_b = array_2_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_18_a = array_2_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_18_valid_a = array_2_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_18_b = array_2_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_19_a = array_2_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_19_valid_a = array_2_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_19_b = array_2_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_20_a = array_2_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_20_valid_a = array_2_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_20_b = array_2_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_21_a = array_2_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_21_valid_a = array_2_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_21_b = array_2_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_22_a = array_2_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_22_valid_a = array_2_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_22_b = array_2_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_23_a = array_2_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_23_valid_a = array_2_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_23_b = array_2_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_24_a = array_2_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_24_valid_a = array_2_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_24_b = array_2_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_25_a = array_2_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_25_valid_a = array_2_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_25_b = array_2_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_26_a = array_2_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_26_valid_a = array_2_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_26_b = array_2_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_27_a = array_2_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_27_valid_a = array_2_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_27_b = array_2_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_28_a = array_2_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_28_valid_a = array_2_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_28_b = array_2_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_29_a = array_2_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_29_valid_a = array_2_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_29_b = array_2_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_30_a = array_2_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_30_valid_a = array_2_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_30_b = array_2_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_3_io_d_in_31_a = array_2_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_31_valid_a = array_2_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_3_io_d_in_31_b = array_2_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_3_io_wr_en_mem1 = io_wr_en_mem1_3; // @[Array.scala 71:28]
  assign array_3_io_wr_en_mem2 = io_wr_en_mem2_3; // @[Array.scala 72:28]
  assign array_3_io_wr_en_mem3 = io_wr_en_mem3_3; // @[Array.scala 73:28]
  assign array_3_io_wr_en_mem4 = io_wr_en_mem4_3; // @[Array.scala 74:28]
  assign array_3_io_wr_en_mem5 = io_wr_en_mem5_3; // @[Array.scala 75:28]
  assign array_3_io_wr_en_mem6 = io_wr_en_mem6_3; // @[Array.scala 76:28]
  assign array_3_io_wr_instr_mem1 = io_wr_instr_mem1_3; // @[Array.scala 77:31]
  assign array_3_io_wr_instr_mem2 = io_wr_instr_mem2_3; // @[Array.scala 78:31]
  assign array_3_io_wr_instr_mem3 = io_wr_instr_mem3_3; // @[Array.scala 79:31]
  assign array_3_io_wr_instr_mem4 = io_wr_instr_mem4_3; // @[Array.scala 80:31]
  assign array_3_io_wr_instr_mem5 = io_wr_instr_mem5_3; // @[Array.scala 81:31]
  assign array_3_io_wr_instr_mem6 = io_wr_instr_mem6_3; // @[Array.scala 82:31]
  assign array_3_io_PC1_in = array_2_io_PC6_out; // @[Array.scala 84:24]
  assign array_3_io_Addr_in = array_2_io_Addr_out; // @[Array.scala 85:25]
  assign array_3_io_Tag_in_Tag = array_2_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_3_io_Tag_in_RoundCnt = array_2_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
  assign array_4_clock = clock;
  assign array_4_reset = reset;
  assign array_4_io_d_in_0_a = array_3_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_0_valid_a = array_3_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_0_b = array_3_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_1_a = array_3_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_1_valid_a = array_3_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_1_b = array_3_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_2_a = array_3_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_2_valid_a = array_3_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_2_b = array_3_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_3_a = array_3_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_3_valid_a = array_3_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_3_b = array_3_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_4_a = array_3_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_4_valid_a = array_3_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_4_b = array_3_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_5_a = array_3_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_5_valid_a = array_3_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_5_b = array_3_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_6_a = array_3_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_6_valid_a = array_3_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_6_b = array_3_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_7_a = array_3_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_7_valid_a = array_3_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_7_b = array_3_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_8_a = array_3_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_8_valid_a = array_3_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_8_b = array_3_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_9_a = array_3_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_9_valid_a = array_3_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_9_b = array_3_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_10_a = array_3_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_10_valid_a = array_3_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_10_b = array_3_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_11_a = array_3_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_11_valid_a = array_3_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_11_b = array_3_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_12_a = array_3_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_12_valid_a = array_3_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_12_b = array_3_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_13_a = array_3_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_13_valid_a = array_3_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_13_b = array_3_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_14_a = array_3_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_14_valid_a = array_3_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_14_b = array_3_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_15_a = array_3_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_15_valid_a = array_3_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_15_b = array_3_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_16_a = array_3_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_16_valid_a = array_3_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_16_b = array_3_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_17_a = array_3_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_17_valid_a = array_3_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_17_b = array_3_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_18_a = array_3_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_18_valid_a = array_3_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_18_b = array_3_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_19_a = array_3_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_19_valid_a = array_3_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_19_b = array_3_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_20_a = array_3_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_20_valid_a = array_3_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_20_b = array_3_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_21_a = array_3_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_21_valid_a = array_3_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_21_b = array_3_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_22_a = array_3_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_22_valid_a = array_3_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_22_b = array_3_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_23_a = array_3_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_23_valid_a = array_3_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_23_b = array_3_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_24_a = array_3_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_24_valid_a = array_3_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_24_b = array_3_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_25_a = array_3_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_25_valid_a = array_3_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_25_b = array_3_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_26_a = array_3_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_26_valid_a = array_3_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_26_b = array_3_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_27_a = array_3_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_27_valid_a = array_3_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_27_b = array_3_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_28_a = array_3_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_28_valid_a = array_3_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_28_b = array_3_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_29_a = array_3_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_29_valid_a = array_3_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_29_b = array_3_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_30_a = array_3_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_30_valid_a = array_3_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_30_b = array_3_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_4_io_d_in_31_a = array_3_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_31_valid_a = array_3_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_4_io_d_in_31_b = array_3_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_4_io_wr_en_mem1 = io_wr_en_mem1_4; // @[Array.scala 71:28]
  assign array_4_io_wr_en_mem2 = io_wr_en_mem2_4; // @[Array.scala 72:28]
  assign array_4_io_wr_en_mem3 = io_wr_en_mem3_4; // @[Array.scala 73:28]
  assign array_4_io_wr_en_mem4 = io_wr_en_mem4_4; // @[Array.scala 74:28]
  assign array_4_io_wr_en_mem5 = io_wr_en_mem5_4; // @[Array.scala 75:28]
  assign array_4_io_wr_en_mem6 = io_wr_en_mem6_4; // @[Array.scala 76:28]
  assign array_4_io_wr_instr_mem1 = io_wr_instr_mem1_4; // @[Array.scala 77:31]
  assign array_4_io_wr_instr_mem2 = io_wr_instr_mem2_4; // @[Array.scala 78:31]
  assign array_4_io_wr_instr_mem3 = io_wr_instr_mem3_4; // @[Array.scala 79:31]
  assign array_4_io_wr_instr_mem4 = io_wr_instr_mem4_4; // @[Array.scala 80:31]
  assign array_4_io_wr_instr_mem5 = io_wr_instr_mem5_4; // @[Array.scala 81:31]
  assign array_4_io_wr_instr_mem6 = io_wr_instr_mem6_4; // @[Array.scala 82:31]
  assign array_4_io_PC1_in = array_3_io_PC6_out; // @[Array.scala 84:24]
  assign array_4_io_Addr_in = array_3_io_Addr_out; // @[Array.scala 85:25]
  assign array_4_io_Tag_in_Tag = array_3_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_4_io_Tag_in_RoundCnt = array_3_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
  assign array_5_clock = clock;
  assign array_5_reset = reset;
  assign array_5_io_d_in_0_a = array_4_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_0_valid_a = array_4_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_0_b = array_4_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_1_a = array_4_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_1_valid_a = array_4_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_1_b = array_4_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_2_a = array_4_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_2_valid_a = array_4_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_2_b = array_4_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_3_a = array_4_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_3_valid_a = array_4_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_3_b = array_4_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_4_a = array_4_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_4_valid_a = array_4_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_4_b = array_4_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_5_a = array_4_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_5_valid_a = array_4_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_5_b = array_4_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_6_a = array_4_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_6_valid_a = array_4_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_6_b = array_4_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_7_a = array_4_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_7_valid_a = array_4_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_7_b = array_4_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_8_a = array_4_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_8_valid_a = array_4_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_8_b = array_4_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_9_a = array_4_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_9_valid_a = array_4_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_9_b = array_4_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_10_a = array_4_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_10_valid_a = array_4_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_10_b = array_4_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_11_a = array_4_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_11_valid_a = array_4_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_11_b = array_4_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_12_a = array_4_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_12_valid_a = array_4_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_12_b = array_4_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_13_a = array_4_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_13_valid_a = array_4_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_13_b = array_4_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_14_a = array_4_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_14_valid_a = array_4_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_14_b = array_4_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_15_a = array_4_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_15_valid_a = array_4_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_15_b = array_4_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_16_a = array_4_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_16_valid_a = array_4_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_16_b = array_4_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_17_a = array_4_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_17_valid_a = array_4_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_17_b = array_4_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_18_a = array_4_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_18_valid_a = array_4_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_18_b = array_4_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_19_a = array_4_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_19_valid_a = array_4_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_19_b = array_4_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_20_a = array_4_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_20_valid_a = array_4_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_20_b = array_4_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_21_a = array_4_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_21_valid_a = array_4_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_21_b = array_4_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_22_a = array_4_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_22_valid_a = array_4_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_22_b = array_4_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_23_a = array_4_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_23_valid_a = array_4_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_23_b = array_4_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_24_a = array_4_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_24_valid_a = array_4_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_24_b = array_4_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_25_a = array_4_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_25_valid_a = array_4_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_25_b = array_4_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_26_a = array_4_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_26_valid_a = array_4_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_26_b = array_4_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_27_a = array_4_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_27_valid_a = array_4_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_27_b = array_4_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_28_a = array_4_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_28_valid_a = array_4_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_28_b = array_4_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_29_a = array_4_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_29_valid_a = array_4_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_29_b = array_4_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_30_a = array_4_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_30_valid_a = array_4_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_30_b = array_4_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_5_io_d_in_31_a = array_4_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_31_valid_a = array_4_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_5_io_d_in_31_b = array_4_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_5_io_wr_en_mem1 = io_wr_en_mem1_5; // @[Array.scala 71:28]
  assign array_5_io_wr_en_mem2 = io_wr_en_mem2_5; // @[Array.scala 72:28]
  assign array_5_io_wr_en_mem3 = io_wr_en_mem3_5; // @[Array.scala 73:28]
  assign array_5_io_wr_en_mem4 = io_wr_en_mem4_5; // @[Array.scala 74:28]
  assign array_5_io_wr_en_mem5 = io_wr_en_mem5_5; // @[Array.scala 75:28]
  assign array_5_io_wr_en_mem6 = io_wr_en_mem6_5; // @[Array.scala 76:28]
  assign array_5_io_wr_instr_mem1 = io_wr_instr_mem1_5; // @[Array.scala 77:31]
  assign array_5_io_wr_instr_mem2 = io_wr_instr_mem2_5; // @[Array.scala 78:31]
  assign array_5_io_wr_instr_mem3 = io_wr_instr_mem3_5; // @[Array.scala 79:31]
  assign array_5_io_wr_instr_mem4 = io_wr_instr_mem4_5; // @[Array.scala 80:31]
  assign array_5_io_wr_instr_mem5 = io_wr_instr_mem5_5; // @[Array.scala 81:31]
  assign array_5_io_wr_instr_mem6 = io_wr_instr_mem6_5; // @[Array.scala 82:31]
  assign array_5_io_PC1_in = array_4_io_PC6_out; // @[Array.scala 84:24]
  assign array_5_io_Addr_in = array_4_io_Addr_out; // @[Array.scala 85:25]
  assign array_5_io_Tag_in_Tag = array_4_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_5_io_Tag_in_RoundCnt = array_4_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
  assign array_6_clock = clock;
  assign array_6_reset = reset;
  assign array_6_io_d_in_0_a = array_5_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_0_valid_a = array_5_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_0_b = array_5_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_1_a = array_5_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_1_valid_a = array_5_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_1_b = array_5_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_2_a = array_5_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_2_valid_a = array_5_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_2_b = array_5_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_3_a = array_5_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_3_valid_a = array_5_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_3_b = array_5_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_4_a = array_5_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_4_valid_a = array_5_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_4_b = array_5_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_5_a = array_5_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_5_valid_a = array_5_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_5_b = array_5_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_6_a = array_5_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_6_valid_a = array_5_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_6_b = array_5_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_7_a = array_5_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_7_valid_a = array_5_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_7_b = array_5_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_8_a = array_5_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_8_valid_a = array_5_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_8_b = array_5_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_9_a = array_5_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_9_valid_a = array_5_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_9_b = array_5_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_10_a = array_5_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_10_valid_a = array_5_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_10_b = array_5_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_11_a = array_5_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_11_valid_a = array_5_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_11_b = array_5_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_12_a = array_5_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_12_valid_a = array_5_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_12_b = array_5_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_13_a = array_5_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_13_valid_a = array_5_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_13_b = array_5_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_14_a = array_5_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_14_valid_a = array_5_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_14_b = array_5_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_15_a = array_5_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_15_valid_a = array_5_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_15_b = array_5_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_16_a = array_5_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_16_valid_a = array_5_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_16_b = array_5_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_17_a = array_5_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_17_valid_a = array_5_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_17_b = array_5_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_18_a = array_5_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_18_valid_a = array_5_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_18_b = array_5_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_19_a = array_5_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_19_valid_a = array_5_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_19_b = array_5_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_20_a = array_5_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_20_valid_a = array_5_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_20_b = array_5_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_21_a = array_5_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_21_valid_a = array_5_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_21_b = array_5_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_22_a = array_5_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_22_valid_a = array_5_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_22_b = array_5_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_23_a = array_5_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_23_valid_a = array_5_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_23_b = array_5_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_24_a = array_5_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_24_valid_a = array_5_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_24_b = array_5_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_25_a = array_5_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_25_valid_a = array_5_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_25_b = array_5_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_26_a = array_5_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_26_valid_a = array_5_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_26_b = array_5_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_27_a = array_5_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_27_valid_a = array_5_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_27_b = array_5_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_28_a = array_5_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_28_valid_a = array_5_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_28_b = array_5_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_29_a = array_5_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_29_valid_a = array_5_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_29_b = array_5_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_30_a = array_5_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_30_valid_a = array_5_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_30_b = array_5_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_6_io_d_in_31_a = array_5_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_31_valid_a = array_5_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_6_io_d_in_31_b = array_5_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_6_io_wr_en_mem1 = io_wr_en_mem1_6; // @[Array.scala 71:28]
  assign array_6_io_wr_en_mem2 = io_wr_en_mem2_6; // @[Array.scala 72:28]
  assign array_6_io_wr_en_mem3 = io_wr_en_mem3_6; // @[Array.scala 73:28]
  assign array_6_io_wr_en_mem4 = io_wr_en_mem4_6; // @[Array.scala 74:28]
  assign array_6_io_wr_en_mem5 = io_wr_en_mem5_6; // @[Array.scala 75:28]
  assign array_6_io_wr_en_mem6 = io_wr_en_mem6_6; // @[Array.scala 76:28]
  assign array_6_io_wr_instr_mem1 = io_wr_instr_mem1_6; // @[Array.scala 77:31]
  assign array_6_io_wr_instr_mem2 = io_wr_instr_mem2_6; // @[Array.scala 78:31]
  assign array_6_io_wr_instr_mem3 = io_wr_instr_mem3_6; // @[Array.scala 79:31]
  assign array_6_io_wr_instr_mem4 = io_wr_instr_mem4_6; // @[Array.scala 80:31]
  assign array_6_io_wr_instr_mem5 = io_wr_instr_mem5_6; // @[Array.scala 81:31]
  assign array_6_io_wr_instr_mem6 = io_wr_instr_mem6_6; // @[Array.scala 82:31]
  assign array_6_io_PC1_in = array_5_io_PC6_out; // @[Array.scala 84:24]
  assign array_6_io_Addr_in = array_5_io_Addr_out; // @[Array.scala 85:25]
  assign array_6_io_Tag_in_Tag = array_5_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_6_io_Tag_in_RoundCnt = array_5_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
  assign array_7_clock = clock;
  assign array_7_reset = reset;
  assign array_7_io_d_in_0_a = array_6_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_0_valid_a = array_6_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_0_b = array_6_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_1_a = array_6_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_1_valid_a = array_6_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_1_b = array_6_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_2_a = array_6_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_2_valid_a = array_6_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_2_b = array_6_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_3_a = array_6_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_3_valid_a = array_6_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_3_b = array_6_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_4_a = array_6_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_4_valid_a = array_6_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_4_b = array_6_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_5_a = array_6_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_5_valid_a = array_6_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_5_b = array_6_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_6_a = array_6_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_6_valid_a = array_6_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_6_b = array_6_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_7_a = array_6_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_7_valid_a = array_6_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_7_b = array_6_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_8_a = array_6_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_8_valid_a = array_6_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_8_b = array_6_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_9_a = array_6_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_9_valid_a = array_6_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_9_b = array_6_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_10_a = array_6_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_10_valid_a = array_6_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_10_b = array_6_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_11_a = array_6_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_11_valid_a = array_6_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_11_b = array_6_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_12_a = array_6_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_12_valid_a = array_6_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_12_b = array_6_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_13_a = array_6_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_13_valid_a = array_6_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_13_b = array_6_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_14_a = array_6_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_14_valid_a = array_6_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_14_b = array_6_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_15_a = array_6_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_15_valid_a = array_6_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_15_b = array_6_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_16_a = array_6_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_16_valid_a = array_6_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_16_b = array_6_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_17_a = array_6_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_17_valid_a = array_6_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_17_b = array_6_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_18_a = array_6_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_18_valid_a = array_6_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_18_b = array_6_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_19_a = array_6_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_19_valid_a = array_6_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_19_b = array_6_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_20_a = array_6_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_20_valid_a = array_6_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_20_b = array_6_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_21_a = array_6_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_21_valid_a = array_6_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_21_b = array_6_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_22_a = array_6_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_22_valid_a = array_6_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_22_b = array_6_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_23_a = array_6_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_23_valid_a = array_6_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_23_b = array_6_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_24_a = array_6_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_24_valid_a = array_6_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_24_b = array_6_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_25_a = array_6_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_25_valid_a = array_6_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_25_b = array_6_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_26_a = array_6_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_26_valid_a = array_6_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_26_b = array_6_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_27_a = array_6_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_27_valid_a = array_6_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_27_b = array_6_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_28_a = array_6_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_28_valid_a = array_6_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_28_b = array_6_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_29_a = array_6_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_29_valid_a = array_6_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_29_b = array_6_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_30_a = array_6_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_30_valid_a = array_6_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_30_b = array_6_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_7_io_d_in_31_a = array_6_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_31_valid_a = array_6_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_7_io_d_in_31_b = array_6_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_7_io_wr_en_mem1 = io_wr_en_mem1_7; // @[Array.scala 71:28]
  assign array_7_io_wr_en_mem2 = io_wr_en_mem2_7; // @[Array.scala 72:28]
  assign array_7_io_wr_en_mem3 = io_wr_en_mem3_7; // @[Array.scala 73:28]
  assign array_7_io_wr_en_mem4 = io_wr_en_mem4_7; // @[Array.scala 74:28]
  assign array_7_io_wr_en_mem5 = io_wr_en_mem5_7; // @[Array.scala 75:28]
  assign array_7_io_wr_en_mem6 = io_wr_en_mem6_7; // @[Array.scala 76:28]
  assign array_7_io_wr_instr_mem1 = io_wr_instr_mem1_7; // @[Array.scala 77:31]
  assign array_7_io_wr_instr_mem2 = io_wr_instr_mem2_7; // @[Array.scala 78:31]
  assign array_7_io_wr_instr_mem3 = io_wr_instr_mem3_7; // @[Array.scala 79:31]
  assign array_7_io_wr_instr_mem4 = io_wr_instr_mem4_7; // @[Array.scala 80:31]
  assign array_7_io_wr_instr_mem5 = io_wr_instr_mem5_7; // @[Array.scala 81:31]
  assign array_7_io_wr_instr_mem6 = io_wr_instr_mem6_7; // @[Array.scala 82:31]
  assign array_7_io_PC1_in = array_6_io_PC6_out; // @[Array.scala 84:24]
  assign array_7_io_Addr_in = array_6_io_Addr_out; // @[Array.scala 85:25]
  assign array_7_io_Tag_in_Tag = array_6_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_7_io_Tag_in_RoundCnt = array_6_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
  assign array_8_clock = clock;
  assign array_8_reset = reset;
  assign array_8_io_d_in_0_a = array_7_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_0_valid_a = array_7_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_0_b = array_7_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_1_a = array_7_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_1_valid_a = array_7_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_1_b = array_7_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_2_a = array_7_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_2_valid_a = array_7_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_2_b = array_7_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_3_a = array_7_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_3_valid_a = array_7_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_3_b = array_7_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_4_a = array_7_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_4_valid_a = array_7_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_4_b = array_7_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_5_a = array_7_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_5_valid_a = array_7_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_5_b = array_7_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_6_a = array_7_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_6_valid_a = array_7_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_6_b = array_7_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_7_a = array_7_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_7_valid_a = array_7_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_7_b = array_7_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_8_a = array_7_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_8_valid_a = array_7_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_8_b = array_7_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_9_a = array_7_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_9_valid_a = array_7_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_9_b = array_7_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_10_a = array_7_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_10_valid_a = array_7_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_10_b = array_7_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_11_a = array_7_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_11_valid_a = array_7_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_11_b = array_7_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_12_a = array_7_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_12_valid_a = array_7_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_12_b = array_7_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_13_a = array_7_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_13_valid_a = array_7_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_13_b = array_7_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_14_a = array_7_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_14_valid_a = array_7_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_14_b = array_7_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_15_a = array_7_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_15_valid_a = array_7_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_15_b = array_7_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_16_a = array_7_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_16_valid_a = array_7_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_16_b = array_7_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_17_a = array_7_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_17_valid_a = array_7_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_17_b = array_7_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_18_a = array_7_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_18_valid_a = array_7_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_18_b = array_7_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_19_a = array_7_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_19_valid_a = array_7_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_19_b = array_7_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_20_a = array_7_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_20_valid_a = array_7_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_20_b = array_7_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_21_a = array_7_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_21_valid_a = array_7_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_21_b = array_7_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_22_a = array_7_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_22_valid_a = array_7_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_22_b = array_7_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_23_a = array_7_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_23_valid_a = array_7_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_23_b = array_7_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_24_a = array_7_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_24_valid_a = array_7_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_24_b = array_7_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_25_a = array_7_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_25_valid_a = array_7_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_25_b = array_7_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_26_a = array_7_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_26_valid_a = array_7_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_26_b = array_7_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_27_a = array_7_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_27_valid_a = array_7_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_27_b = array_7_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_28_a = array_7_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_28_valid_a = array_7_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_28_b = array_7_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_29_a = array_7_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_29_valid_a = array_7_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_29_b = array_7_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_30_a = array_7_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_30_valid_a = array_7_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_30_b = array_7_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_8_io_d_in_31_a = array_7_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_31_valid_a = array_7_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_8_io_d_in_31_b = array_7_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_8_io_wr_en_mem1 = io_wr_en_mem1_8; // @[Array.scala 71:28]
  assign array_8_io_wr_en_mem2 = io_wr_en_mem2_8; // @[Array.scala 72:28]
  assign array_8_io_wr_en_mem3 = io_wr_en_mem3_8; // @[Array.scala 73:28]
  assign array_8_io_wr_en_mem4 = io_wr_en_mem4_8; // @[Array.scala 74:28]
  assign array_8_io_wr_en_mem5 = io_wr_en_mem5_8; // @[Array.scala 75:28]
  assign array_8_io_wr_en_mem6 = io_wr_en_mem6_8; // @[Array.scala 76:28]
  assign array_8_io_wr_instr_mem1 = io_wr_instr_mem1_8; // @[Array.scala 77:31]
  assign array_8_io_wr_instr_mem2 = io_wr_instr_mem2_8; // @[Array.scala 78:31]
  assign array_8_io_wr_instr_mem3 = io_wr_instr_mem3_8; // @[Array.scala 79:31]
  assign array_8_io_wr_instr_mem4 = io_wr_instr_mem4_8; // @[Array.scala 80:31]
  assign array_8_io_wr_instr_mem5 = io_wr_instr_mem5_8; // @[Array.scala 81:31]
  assign array_8_io_wr_instr_mem6 = io_wr_instr_mem6_8; // @[Array.scala 82:31]
  assign array_8_io_PC1_in = array_7_io_PC6_out; // @[Array.scala 84:24]
  assign array_8_io_Addr_in = array_7_io_Addr_out; // @[Array.scala 85:25]
  assign array_8_io_Tag_in_Tag = array_7_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_8_io_Tag_in_RoundCnt = array_7_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
  assign array_9_clock = clock;
  assign array_9_reset = reset;
  assign array_9_io_d_in_0_a = array_8_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_0_valid_a = array_8_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_0_b = array_8_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_1_a = array_8_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_1_valid_a = array_8_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_1_b = array_8_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_2_a = array_8_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_2_valid_a = array_8_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_2_b = array_8_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_3_a = array_8_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_3_valid_a = array_8_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_3_b = array_8_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_4_a = array_8_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_4_valid_a = array_8_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_4_b = array_8_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_5_a = array_8_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_5_valid_a = array_8_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_5_b = array_8_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_6_a = array_8_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_6_valid_a = array_8_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_6_b = array_8_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_7_a = array_8_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_7_valid_a = array_8_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_7_b = array_8_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_8_a = array_8_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_8_valid_a = array_8_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_8_b = array_8_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_9_a = array_8_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_9_valid_a = array_8_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_9_b = array_8_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_10_a = array_8_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_10_valid_a = array_8_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_10_b = array_8_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_11_a = array_8_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_11_valid_a = array_8_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_11_b = array_8_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_12_a = array_8_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_12_valid_a = array_8_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_12_b = array_8_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_13_a = array_8_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_13_valid_a = array_8_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_13_b = array_8_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_14_a = array_8_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_14_valid_a = array_8_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_14_b = array_8_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_15_a = array_8_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_15_valid_a = array_8_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_15_b = array_8_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_16_a = array_8_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_16_valid_a = array_8_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_16_b = array_8_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_17_a = array_8_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_17_valid_a = array_8_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_17_b = array_8_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_18_a = array_8_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_18_valid_a = array_8_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_18_b = array_8_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_19_a = array_8_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_19_valid_a = array_8_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_19_b = array_8_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_20_a = array_8_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_20_valid_a = array_8_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_20_b = array_8_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_21_a = array_8_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_21_valid_a = array_8_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_21_b = array_8_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_22_a = array_8_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_22_valid_a = array_8_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_22_b = array_8_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_23_a = array_8_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_23_valid_a = array_8_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_23_b = array_8_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_24_a = array_8_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_24_valid_a = array_8_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_24_b = array_8_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_25_a = array_8_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_25_valid_a = array_8_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_25_b = array_8_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_26_a = array_8_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_26_valid_a = array_8_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_26_b = array_8_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_27_a = array_8_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_27_valid_a = array_8_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_27_b = array_8_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_28_a = array_8_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_28_valid_a = array_8_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_28_b = array_8_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_29_a = array_8_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_29_valid_a = array_8_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_29_b = array_8_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_30_a = array_8_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_30_valid_a = array_8_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_30_b = array_8_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_9_io_d_in_31_a = array_8_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_31_valid_a = array_8_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_9_io_d_in_31_b = array_8_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_9_io_wr_en_mem1 = io_wr_en_mem1_9; // @[Array.scala 71:28]
  assign array_9_io_wr_en_mem2 = io_wr_en_mem2_9; // @[Array.scala 72:28]
  assign array_9_io_wr_en_mem3 = io_wr_en_mem3_9; // @[Array.scala 73:28]
  assign array_9_io_wr_en_mem4 = io_wr_en_mem4_9; // @[Array.scala 74:28]
  assign array_9_io_wr_en_mem5 = io_wr_en_mem5_9; // @[Array.scala 75:28]
  assign array_9_io_wr_en_mem6 = io_wr_en_mem6_9; // @[Array.scala 76:28]
  assign array_9_io_wr_instr_mem1 = io_wr_instr_mem1_9; // @[Array.scala 77:31]
  assign array_9_io_wr_instr_mem2 = io_wr_instr_mem2_9; // @[Array.scala 78:31]
  assign array_9_io_wr_instr_mem3 = io_wr_instr_mem3_9; // @[Array.scala 79:31]
  assign array_9_io_wr_instr_mem4 = io_wr_instr_mem4_9; // @[Array.scala 80:31]
  assign array_9_io_wr_instr_mem5 = io_wr_instr_mem5_9; // @[Array.scala 81:31]
  assign array_9_io_wr_instr_mem6 = io_wr_instr_mem6_9; // @[Array.scala 82:31]
  assign array_9_io_PC1_in = array_8_io_PC6_out; // @[Array.scala 84:24]
  assign array_9_io_Addr_in = array_8_io_Addr_out; // @[Array.scala 85:25]
  assign array_9_io_Tag_in_Tag = array_8_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_9_io_Tag_in_RoundCnt = array_8_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
  assign array_10_clock = clock;
  assign array_10_reset = reset;
  assign array_10_io_d_in_0_a = array_9_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_0_valid_a = array_9_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_0_b = array_9_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_1_a = array_9_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_1_valid_a = array_9_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_1_b = array_9_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_2_a = array_9_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_2_valid_a = array_9_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_2_b = array_9_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_3_a = array_9_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_3_valid_a = array_9_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_3_b = array_9_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_4_a = array_9_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_4_valid_a = array_9_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_4_b = array_9_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_5_a = array_9_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_5_valid_a = array_9_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_5_b = array_9_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_6_a = array_9_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_6_valid_a = array_9_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_6_b = array_9_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_7_a = array_9_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_7_valid_a = array_9_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_7_b = array_9_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_8_a = array_9_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_8_valid_a = array_9_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_8_b = array_9_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_9_a = array_9_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_9_valid_a = array_9_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_9_b = array_9_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_10_a = array_9_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_10_valid_a = array_9_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_10_b = array_9_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_11_a = array_9_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_11_valid_a = array_9_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_11_b = array_9_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_12_a = array_9_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_12_valid_a = array_9_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_12_b = array_9_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_13_a = array_9_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_13_valid_a = array_9_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_13_b = array_9_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_14_a = array_9_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_14_valid_a = array_9_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_14_b = array_9_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_15_a = array_9_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_15_valid_a = array_9_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_15_b = array_9_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_16_a = array_9_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_16_valid_a = array_9_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_16_b = array_9_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_17_a = array_9_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_17_valid_a = array_9_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_17_b = array_9_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_18_a = array_9_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_18_valid_a = array_9_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_18_b = array_9_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_19_a = array_9_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_19_valid_a = array_9_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_19_b = array_9_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_20_a = array_9_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_20_valid_a = array_9_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_20_b = array_9_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_21_a = array_9_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_21_valid_a = array_9_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_21_b = array_9_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_22_a = array_9_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_22_valid_a = array_9_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_22_b = array_9_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_23_a = array_9_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_23_valid_a = array_9_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_23_b = array_9_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_24_a = array_9_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_24_valid_a = array_9_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_24_b = array_9_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_25_a = array_9_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_25_valid_a = array_9_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_25_b = array_9_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_26_a = array_9_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_26_valid_a = array_9_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_26_b = array_9_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_27_a = array_9_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_27_valid_a = array_9_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_27_b = array_9_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_28_a = array_9_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_28_valid_a = array_9_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_28_b = array_9_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_29_a = array_9_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_29_valid_a = array_9_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_29_b = array_9_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_30_a = array_9_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_30_valid_a = array_9_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_30_b = array_9_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_10_io_d_in_31_a = array_9_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_31_valid_a = array_9_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_10_io_d_in_31_b = array_9_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_10_io_wr_en_mem1 = io_wr_en_mem1_10; // @[Array.scala 71:28]
  assign array_10_io_wr_en_mem2 = io_wr_en_mem2_10; // @[Array.scala 72:28]
  assign array_10_io_wr_en_mem3 = io_wr_en_mem3_10; // @[Array.scala 73:28]
  assign array_10_io_wr_en_mem4 = io_wr_en_mem4_10; // @[Array.scala 74:28]
  assign array_10_io_wr_en_mem5 = io_wr_en_mem5_10; // @[Array.scala 75:28]
  assign array_10_io_wr_en_mem6 = io_wr_en_mem6_10; // @[Array.scala 76:28]
  assign array_10_io_wr_instr_mem1 = io_wr_instr_mem1_10; // @[Array.scala 77:31]
  assign array_10_io_wr_instr_mem2 = io_wr_instr_mem2_10; // @[Array.scala 78:31]
  assign array_10_io_wr_instr_mem3 = io_wr_instr_mem3_10; // @[Array.scala 79:31]
  assign array_10_io_wr_instr_mem4 = io_wr_instr_mem4_10; // @[Array.scala 80:31]
  assign array_10_io_wr_instr_mem5 = io_wr_instr_mem5_10; // @[Array.scala 81:31]
  assign array_10_io_wr_instr_mem6 = io_wr_instr_mem6_10; // @[Array.scala 82:31]
  assign array_10_io_PC1_in = array_9_io_PC6_out; // @[Array.scala 84:24]
  assign array_10_io_Addr_in = array_9_io_Addr_out; // @[Array.scala 85:25]
  assign array_10_io_Tag_in_Tag = array_9_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_10_io_Tag_in_RoundCnt = array_9_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
  assign array_11_clock = clock;
  assign array_11_reset = reset;
  assign array_11_io_d_in_0_a = array_10_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_0_valid_a = array_10_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_0_b = array_10_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_1_a = array_10_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_1_valid_a = array_10_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_1_b = array_10_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_2_a = array_10_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_2_valid_a = array_10_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_2_b = array_10_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_3_a = array_10_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_3_valid_a = array_10_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_3_b = array_10_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_4_a = array_10_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_4_valid_a = array_10_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_4_b = array_10_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_5_a = array_10_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_5_valid_a = array_10_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_5_b = array_10_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_6_a = array_10_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_6_valid_a = array_10_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_6_b = array_10_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_7_a = array_10_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_7_valid_a = array_10_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_7_b = array_10_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_8_a = array_10_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_8_valid_a = array_10_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_8_b = array_10_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_9_a = array_10_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_9_valid_a = array_10_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_9_b = array_10_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_10_a = array_10_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_10_valid_a = array_10_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_10_b = array_10_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_11_a = array_10_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_11_valid_a = array_10_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_11_b = array_10_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_12_a = array_10_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_12_valid_a = array_10_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_12_b = array_10_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_13_a = array_10_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_13_valid_a = array_10_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_13_b = array_10_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_14_a = array_10_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_14_valid_a = array_10_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_14_b = array_10_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_15_a = array_10_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_15_valid_a = array_10_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_15_b = array_10_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_16_a = array_10_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_16_valid_a = array_10_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_16_b = array_10_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_17_a = array_10_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_17_valid_a = array_10_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_17_b = array_10_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_18_a = array_10_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_18_valid_a = array_10_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_18_b = array_10_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_19_a = array_10_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_19_valid_a = array_10_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_19_b = array_10_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_20_a = array_10_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_20_valid_a = array_10_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_20_b = array_10_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_21_a = array_10_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_21_valid_a = array_10_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_21_b = array_10_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_22_a = array_10_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_22_valid_a = array_10_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_22_b = array_10_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_23_a = array_10_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_23_valid_a = array_10_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_23_b = array_10_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_24_a = array_10_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_24_valid_a = array_10_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_24_b = array_10_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_25_a = array_10_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_25_valid_a = array_10_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_25_b = array_10_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_26_a = array_10_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_26_valid_a = array_10_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_26_b = array_10_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_27_a = array_10_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_27_valid_a = array_10_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_27_b = array_10_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_28_a = array_10_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_28_valid_a = array_10_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_28_b = array_10_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_29_a = array_10_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_29_valid_a = array_10_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_29_b = array_10_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_30_a = array_10_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_30_valid_a = array_10_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_30_b = array_10_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_11_io_d_in_31_a = array_10_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_31_valid_a = array_10_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_11_io_d_in_31_b = array_10_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_11_io_wr_en_mem1 = io_wr_en_mem1_11; // @[Array.scala 71:28]
  assign array_11_io_wr_en_mem2 = io_wr_en_mem2_11; // @[Array.scala 72:28]
  assign array_11_io_wr_en_mem3 = io_wr_en_mem3_11; // @[Array.scala 73:28]
  assign array_11_io_wr_en_mem4 = io_wr_en_mem4_11; // @[Array.scala 74:28]
  assign array_11_io_wr_en_mem5 = io_wr_en_mem5_11; // @[Array.scala 75:28]
  assign array_11_io_wr_en_mem6 = io_wr_en_mem6_11; // @[Array.scala 76:28]
  assign array_11_io_wr_instr_mem1 = io_wr_instr_mem1_11; // @[Array.scala 77:31]
  assign array_11_io_wr_instr_mem2 = io_wr_instr_mem2_11; // @[Array.scala 78:31]
  assign array_11_io_wr_instr_mem3 = io_wr_instr_mem3_11; // @[Array.scala 79:31]
  assign array_11_io_wr_instr_mem4 = io_wr_instr_mem4_11; // @[Array.scala 80:31]
  assign array_11_io_wr_instr_mem5 = io_wr_instr_mem5_11; // @[Array.scala 81:31]
  assign array_11_io_wr_instr_mem6 = io_wr_instr_mem6_11; // @[Array.scala 82:31]
  assign array_11_io_PC1_in = array_10_io_PC6_out; // @[Array.scala 84:24]
  assign array_11_io_Addr_in = array_10_io_Addr_out; // @[Array.scala 85:25]
  assign array_11_io_Tag_in_Tag = array_10_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_11_io_Tag_in_RoundCnt = array_10_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
  assign array_12_clock = clock;
  assign array_12_reset = reset;
  assign array_12_io_d_in_0_a = array_11_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_0_valid_a = array_11_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_0_b = array_11_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_1_a = array_11_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_1_valid_a = array_11_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_1_b = array_11_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_2_a = array_11_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_2_valid_a = array_11_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_2_b = array_11_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_3_a = array_11_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_3_valid_a = array_11_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_3_b = array_11_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_4_a = array_11_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_4_valid_a = array_11_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_4_b = array_11_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_5_a = array_11_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_5_valid_a = array_11_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_5_b = array_11_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_6_a = array_11_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_6_valid_a = array_11_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_6_b = array_11_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_7_a = array_11_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_7_valid_a = array_11_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_7_b = array_11_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_8_a = array_11_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_8_valid_a = array_11_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_8_b = array_11_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_9_a = array_11_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_9_valid_a = array_11_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_9_b = array_11_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_10_a = array_11_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_10_valid_a = array_11_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_10_b = array_11_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_11_a = array_11_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_11_valid_a = array_11_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_11_b = array_11_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_12_a = array_11_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_12_valid_a = array_11_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_12_b = array_11_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_13_a = array_11_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_13_valid_a = array_11_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_13_b = array_11_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_14_a = array_11_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_14_valid_a = array_11_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_14_b = array_11_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_15_a = array_11_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_15_valid_a = array_11_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_15_b = array_11_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_16_a = array_11_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_16_valid_a = array_11_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_16_b = array_11_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_17_a = array_11_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_17_valid_a = array_11_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_17_b = array_11_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_18_a = array_11_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_18_valid_a = array_11_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_18_b = array_11_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_19_a = array_11_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_19_valid_a = array_11_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_19_b = array_11_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_20_a = array_11_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_20_valid_a = array_11_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_20_b = array_11_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_21_a = array_11_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_21_valid_a = array_11_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_21_b = array_11_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_22_a = array_11_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_22_valid_a = array_11_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_22_b = array_11_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_23_a = array_11_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_23_valid_a = array_11_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_23_b = array_11_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_24_a = array_11_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_24_valid_a = array_11_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_24_b = array_11_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_25_a = array_11_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_25_valid_a = array_11_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_25_b = array_11_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_26_a = array_11_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_26_valid_a = array_11_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_26_b = array_11_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_27_a = array_11_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_27_valid_a = array_11_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_27_b = array_11_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_28_a = array_11_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_28_valid_a = array_11_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_28_b = array_11_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_29_a = array_11_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_29_valid_a = array_11_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_29_b = array_11_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_30_a = array_11_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_30_valid_a = array_11_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_30_b = array_11_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_12_io_d_in_31_a = array_11_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_31_valid_a = array_11_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_12_io_d_in_31_b = array_11_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_12_io_wr_en_mem1 = io_wr_en_mem1_12; // @[Array.scala 71:28]
  assign array_12_io_wr_en_mem2 = io_wr_en_mem2_12; // @[Array.scala 72:28]
  assign array_12_io_wr_en_mem3 = io_wr_en_mem3_12; // @[Array.scala 73:28]
  assign array_12_io_wr_en_mem4 = io_wr_en_mem4_12; // @[Array.scala 74:28]
  assign array_12_io_wr_en_mem5 = io_wr_en_mem5_12; // @[Array.scala 75:28]
  assign array_12_io_wr_en_mem6 = io_wr_en_mem6_12; // @[Array.scala 76:28]
  assign array_12_io_wr_instr_mem1 = io_wr_instr_mem1_12; // @[Array.scala 77:31]
  assign array_12_io_wr_instr_mem2 = io_wr_instr_mem2_12; // @[Array.scala 78:31]
  assign array_12_io_wr_instr_mem3 = io_wr_instr_mem3_12; // @[Array.scala 79:31]
  assign array_12_io_wr_instr_mem4 = io_wr_instr_mem4_12; // @[Array.scala 80:31]
  assign array_12_io_wr_instr_mem5 = io_wr_instr_mem5_12; // @[Array.scala 81:31]
  assign array_12_io_wr_instr_mem6 = io_wr_instr_mem6_12; // @[Array.scala 82:31]
  assign array_12_io_PC1_in = array_11_io_PC6_out; // @[Array.scala 84:24]
  assign array_12_io_Addr_in = array_11_io_Addr_out; // @[Array.scala 85:25]
  assign array_12_io_Tag_in_Tag = array_11_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_12_io_Tag_in_RoundCnt = array_11_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
  assign array_13_clock = clock;
  assign array_13_reset = reset;
  assign array_13_io_d_in_0_a = array_12_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_0_valid_a = array_12_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_0_b = array_12_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_1_a = array_12_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_1_valid_a = array_12_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_1_b = array_12_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_2_a = array_12_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_2_valid_a = array_12_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_2_b = array_12_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_3_a = array_12_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_3_valid_a = array_12_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_3_b = array_12_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_4_a = array_12_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_4_valid_a = array_12_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_4_b = array_12_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_5_a = array_12_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_5_valid_a = array_12_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_5_b = array_12_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_6_a = array_12_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_6_valid_a = array_12_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_6_b = array_12_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_7_a = array_12_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_7_valid_a = array_12_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_7_b = array_12_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_8_a = array_12_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_8_valid_a = array_12_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_8_b = array_12_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_9_a = array_12_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_9_valid_a = array_12_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_9_b = array_12_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_10_a = array_12_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_10_valid_a = array_12_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_10_b = array_12_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_11_a = array_12_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_11_valid_a = array_12_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_11_b = array_12_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_12_a = array_12_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_12_valid_a = array_12_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_12_b = array_12_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_13_a = array_12_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_13_valid_a = array_12_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_13_b = array_12_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_14_a = array_12_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_14_valid_a = array_12_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_14_b = array_12_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_15_a = array_12_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_15_valid_a = array_12_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_15_b = array_12_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_16_a = array_12_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_16_valid_a = array_12_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_16_b = array_12_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_17_a = array_12_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_17_valid_a = array_12_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_17_b = array_12_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_18_a = array_12_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_18_valid_a = array_12_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_18_b = array_12_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_19_a = array_12_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_19_valid_a = array_12_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_19_b = array_12_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_20_a = array_12_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_20_valid_a = array_12_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_20_b = array_12_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_21_a = array_12_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_21_valid_a = array_12_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_21_b = array_12_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_22_a = array_12_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_22_valid_a = array_12_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_22_b = array_12_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_23_a = array_12_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_23_valid_a = array_12_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_23_b = array_12_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_24_a = array_12_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_24_valid_a = array_12_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_24_b = array_12_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_25_a = array_12_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_25_valid_a = array_12_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_25_b = array_12_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_26_a = array_12_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_26_valid_a = array_12_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_26_b = array_12_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_27_a = array_12_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_27_valid_a = array_12_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_27_b = array_12_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_28_a = array_12_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_28_valid_a = array_12_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_28_b = array_12_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_29_a = array_12_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_29_valid_a = array_12_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_29_b = array_12_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_30_a = array_12_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_30_valid_a = array_12_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_30_b = array_12_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_13_io_d_in_31_a = array_12_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_31_valid_a = array_12_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_13_io_d_in_31_b = array_12_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_13_io_wr_en_mem1 = io_wr_en_mem1_13; // @[Array.scala 71:28]
  assign array_13_io_wr_en_mem2 = io_wr_en_mem2_13; // @[Array.scala 72:28]
  assign array_13_io_wr_en_mem3 = io_wr_en_mem3_13; // @[Array.scala 73:28]
  assign array_13_io_wr_en_mem4 = io_wr_en_mem4_13; // @[Array.scala 74:28]
  assign array_13_io_wr_en_mem5 = io_wr_en_mem5_13; // @[Array.scala 75:28]
  assign array_13_io_wr_en_mem6 = io_wr_en_mem6_13; // @[Array.scala 76:28]
  assign array_13_io_wr_instr_mem1 = io_wr_instr_mem1_13; // @[Array.scala 77:31]
  assign array_13_io_wr_instr_mem2 = io_wr_instr_mem2_13; // @[Array.scala 78:31]
  assign array_13_io_wr_instr_mem3 = io_wr_instr_mem3_13; // @[Array.scala 79:31]
  assign array_13_io_wr_instr_mem4 = io_wr_instr_mem4_13; // @[Array.scala 80:31]
  assign array_13_io_wr_instr_mem5 = io_wr_instr_mem5_13; // @[Array.scala 81:31]
  assign array_13_io_wr_instr_mem6 = io_wr_instr_mem6_13; // @[Array.scala 82:31]
  assign array_13_io_PC1_in = array_12_io_PC6_out; // @[Array.scala 84:24]
  assign array_13_io_Addr_in = array_12_io_Addr_out; // @[Array.scala 85:25]
  assign array_13_io_Tag_in_Tag = array_12_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_13_io_Tag_in_RoundCnt = array_12_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
  assign array_14_clock = clock;
  assign array_14_reset = reset;
  assign array_14_io_d_in_0_a = array_13_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_0_valid_a = array_13_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_0_b = array_13_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_1_a = array_13_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_1_valid_a = array_13_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_1_b = array_13_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_2_a = array_13_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_2_valid_a = array_13_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_2_b = array_13_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_3_a = array_13_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_3_valid_a = array_13_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_3_b = array_13_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_4_a = array_13_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_4_valid_a = array_13_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_4_b = array_13_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_5_a = array_13_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_5_valid_a = array_13_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_5_b = array_13_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_6_a = array_13_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_6_valid_a = array_13_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_6_b = array_13_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_7_a = array_13_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_7_valid_a = array_13_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_7_b = array_13_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_8_a = array_13_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_8_valid_a = array_13_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_8_b = array_13_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_9_a = array_13_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_9_valid_a = array_13_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_9_b = array_13_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_10_a = array_13_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_10_valid_a = array_13_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_10_b = array_13_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_11_a = array_13_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_11_valid_a = array_13_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_11_b = array_13_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_12_a = array_13_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_12_valid_a = array_13_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_12_b = array_13_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_13_a = array_13_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_13_valid_a = array_13_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_13_b = array_13_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_14_a = array_13_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_14_valid_a = array_13_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_14_b = array_13_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_15_a = array_13_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_15_valid_a = array_13_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_15_b = array_13_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_16_a = array_13_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_16_valid_a = array_13_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_16_b = array_13_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_17_a = array_13_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_17_valid_a = array_13_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_17_b = array_13_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_18_a = array_13_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_18_valid_a = array_13_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_18_b = array_13_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_19_a = array_13_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_19_valid_a = array_13_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_19_b = array_13_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_20_a = array_13_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_20_valid_a = array_13_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_20_b = array_13_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_21_a = array_13_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_21_valid_a = array_13_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_21_b = array_13_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_22_a = array_13_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_22_valid_a = array_13_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_22_b = array_13_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_23_a = array_13_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_23_valid_a = array_13_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_23_b = array_13_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_24_a = array_13_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_24_valid_a = array_13_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_24_b = array_13_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_25_a = array_13_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_25_valid_a = array_13_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_25_b = array_13_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_26_a = array_13_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_26_valid_a = array_13_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_26_b = array_13_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_27_a = array_13_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_27_valid_a = array_13_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_27_b = array_13_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_28_a = array_13_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_28_valid_a = array_13_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_28_b = array_13_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_29_a = array_13_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_29_valid_a = array_13_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_29_b = array_13_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_30_a = array_13_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_30_valid_a = array_13_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_30_b = array_13_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_14_io_d_in_31_a = array_13_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_31_valid_a = array_13_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_14_io_d_in_31_b = array_13_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_14_io_wr_en_mem1 = io_wr_en_mem1_14; // @[Array.scala 71:28]
  assign array_14_io_wr_en_mem2 = io_wr_en_mem2_14; // @[Array.scala 72:28]
  assign array_14_io_wr_en_mem3 = io_wr_en_mem3_14; // @[Array.scala 73:28]
  assign array_14_io_wr_en_mem4 = io_wr_en_mem4_14; // @[Array.scala 74:28]
  assign array_14_io_wr_en_mem5 = io_wr_en_mem5_14; // @[Array.scala 75:28]
  assign array_14_io_wr_en_mem6 = io_wr_en_mem6_14; // @[Array.scala 76:28]
  assign array_14_io_wr_instr_mem1 = io_wr_instr_mem1_14; // @[Array.scala 77:31]
  assign array_14_io_wr_instr_mem2 = io_wr_instr_mem2_14; // @[Array.scala 78:31]
  assign array_14_io_wr_instr_mem3 = io_wr_instr_mem3_14; // @[Array.scala 79:31]
  assign array_14_io_wr_instr_mem4 = io_wr_instr_mem4_14; // @[Array.scala 80:31]
  assign array_14_io_wr_instr_mem5 = io_wr_instr_mem5_14; // @[Array.scala 81:31]
  assign array_14_io_wr_instr_mem6 = io_wr_instr_mem6_14; // @[Array.scala 82:31]
  assign array_14_io_PC1_in = array_13_io_PC6_out; // @[Array.scala 84:24]
  assign array_14_io_Addr_in = array_13_io_Addr_out; // @[Array.scala 85:25]
  assign array_14_io_Tag_in_Tag = array_13_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_14_io_Tag_in_RoundCnt = array_13_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
  assign array_15_clock = clock;
  assign array_15_reset = reset;
  assign array_15_io_d_in_0_a = array_14_io_d_out_0_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_0_valid_a = array_14_io_d_out_0_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_0_b = array_14_io_d_out_0_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_1_a = array_14_io_d_out_1_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_1_valid_a = array_14_io_d_out_1_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_1_b = array_14_io_d_out_1_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_2_a = array_14_io_d_out_2_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_2_valid_a = array_14_io_d_out_2_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_2_b = array_14_io_d_out_2_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_3_a = array_14_io_d_out_3_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_3_valid_a = array_14_io_d_out_3_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_3_b = array_14_io_d_out_3_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_4_a = array_14_io_d_out_4_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_4_valid_a = array_14_io_d_out_4_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_4_b = array_14_io_d_out_4_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_5_a = array_14_io_d_out_5_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_5_valid_a = array_14_io_d_out_5_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_5_b = array_14_io_d_out_5_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_6_a = array_14_io_d_out_6_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_6_valid_a = array_14_io_d_out_6_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_6_b = array_14_io_d_out_6_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_7_a = array_14_io_d_out_7_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_7_valid_a = array_14_io_d_out_7_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_7_b = array_14_io_d_out_7_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_8_a = array_14_io_d_out_8_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_8_valid_a = array_14_io_d_out_8_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_8_b = array_14_io_d_out_8_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_9_a = array_14_io_d_out_9_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_9_valid_a = array_14_io_d_out_9_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_9_b = array_14_io_d_out_9_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_10_a = array_14_io_d_out_10_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_10_valid_a = array_14_io_d_out_10_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_10_b = array_14_io_d_out_10_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_11_a = array_14_io_d_out_11_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_11_valid_a = array_14_io_d_out_11_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_11_b = array_14_io_d_out_11_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_12_a = array_14_io_d_out_12_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_12_valid_a = array_14_io_d_out_12_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_12_b = array_14_io_d_out_12_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_13_a = array_14_io_d_out_13_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_13_valid_a = array_14_io_d_out_13_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_13_b = array_14_io_d_out_13_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_14_a = array_14_io_d_out_14_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_14_valid_a = array_14_io_d_out_14_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_14_b = array_14_io_d_out_14_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_15_a = array_14_io_d_out_15_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_15_valid_a = array_14_io_d_out_15_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_15_b = array_14_io_d_out_15_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_16_a = array_14_io_d_out_16_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_16_valid_a = array_14_io_d_out_16_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_16_b = array_14_io_d_out_16_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_17_a = array_14_io_d_out_17_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_17_valid_a = array_14_io_d_out_17_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_17_b = array_14_io_d_out_17_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_18_a = array_14_io_d_out_18_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_18_valid_a = array_14_io_d_out_18_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_18_b = array_14_io_d_out_18_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_19_a = array_14_io_d_out_19_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_19_valid_a = array_14_io_d_out_19_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_19_b = array_14_io_d_out_19_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_20_a = array_14_io_d_out_20_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_20_valid_a = array_14_io_d_out_20_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_20_b = array_14_io_d_out_20_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_21_a = array_14_io_d_out_21_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_21_valid_a = array_14_io_d_out_21_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_21_b = array_14_io_d_out_21_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_22_a = array_14_io_d_out_22_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_22_valid_a = array_14_io_d_out_22_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_22_b = array_14_io_d_out_22_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_23_a = array_14_io_d_out_23_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_23_valid_a = array_14_io_d_out_23_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_23_b = array_14_io_d_out_23_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_24_a = array_14_io_d_out_24_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_24_valid_a = array_14_io_d_out_24_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_24_b = array_14_io_d_out_24_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_25_a = array_14_io_d_out_25_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_25_valid_a = array_14_io_d_out_25_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_25_b = array_14_io_d_out_25_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_26_a = array_14_io_d_out_26_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_26_valid_a = array_14_io_d_out_26_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_26_b = array_14_io_d_out_26_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_27_a = array_14_io_d_out_27_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_27_valid_a = array_14_io_d_out_27_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_27_b = array_14_io_d_out_27_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_28_a = array_14_io_d_out_28_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_28_valid_a = array_14_io_d_out_28_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_28_b = array_14_io_d_out_28_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_29_a = array_14_io_d_out_29_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_29_valid_a = array_14_io_d_out_29_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_29_b = array_14_io_d_out_29_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_30_a = array_14_io_d_out_30_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_30_valid_a = array_14_io_d_out_30_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_30_b = array_14_io_d_out_30_b; // @[Array.scala 69:22]
  assign array_15_io_d_in_31_a = array_14_io_d_out_31_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_31_valid_a = array_14_io_d_out_31_valid_a; // @[Array.scala 69:22]
  assign array_15_io_d_in_31_b = array_14_io_d_out_31_b; // @[Array.scala 69:22]
  assign array_15_io_wr_en_mem1 = io_wr_en_mem1_15; // @[Array.scala 71:28]
  assign array_15_io_wr_en_mem2 = io_wr_en_mem2_15; // @[Array.scala 72:28]
  assign array_15_io_wr_en_mem3 = io_wr_en_mem3_15; // @[Array.scala 73:28]
  assign array_15_io_wr_en_mem4 = io_wr_en_mem4_15; // @[Array.scala 74:28]
  assign array_15_io_wr_en_mem5 = io_wr_en_mem5_15; // @[Array.scala 75:28]
  assign array_15_io_wr_en_mem6 = io_wr_en_mem6_15; // @[Array.scala 76:28]
  assign array_15_io_wr_instr_mem1 = io_wr_instr_mem1_15; // @[Array.scala 77:31]
  assign array_15_io_wr_instr_mem2 = io_wr_instr_mem2_15; // @[Array.scala 78:31]
  assign array_15_io_wr_instr_mem3 = io_wr_instr_mem3_15; // @[Array.scala 79:31]
  assign array_15_io_wr_instr_mem4 = io_wr_instr_mem4_15; // @[Array.scala 80:31]
  assign array_15_io_wr_instr_mem5 = io_wr_instr_mem5_15; // @[Array.scala 81:31]
  assign array_15_io_wr_instr_mem6 = io_wr_instr_mem6_15; // @[Array.scala 82:31]
  assign array_15_io_PC1_in = array_14_io_PC6_out; // @[Array.scala 84:24]
  assign array_15_io_Addr_in = array_14_io_Addr_out; // @[Array.scala 85:25]
  assign array_15_io_Tag_in_Tag = array_14_io_Tag_out_Tag; // @[Array.scala 70:24]
  assign array_15_io_Tag_in_RoundCnt = array_14_io_Tag_out_RoundCnt; // @[Array.scala 70:24]
endmodule
module Mem1(
  input  [7:0]   R0_addr,
  input          R0_clk,
  output [287:0] R0_data,
  input  [7:0]   W0_addr,
  input          W0_en,
  input          W0_clk,
  input  [287:0] W0_data
);
  wire [7:0] Mem1_ext_R0_addr;
  wire  Mem1_ext_R0_en;
  wire  Mem1_ext_R0_clk;
  wire [287:0] Mem1_ext_R0_data;
  wire [7:0] Mem1_ext_W0_addr;
  wire  Mem1_ext_W0_en;
  wire  Mem1_ext_W0_clk;
  wire [287:0] Mem1_ext_W0_data;
  Mem1_ext Mem1_ext (
    .R0_addr(Mem1_ext_R0_addr),
    .R0_en(Mem1_ext_R0_en),
    .R0_clk(Mem1_ext_R0_clk),
    .R0_data(Mem1_ext_R0_data),
    .W0_addr(Mem1_ext_W0_addr),
    .W0_en(Mem1_ext_W0_en),
    .W0_clk(Mem1_ext_W0_clk),
    .W0_data(Mem1_ext_W0_data)
  );
  assign Mem1_ext_R0_clk = R0_clk;
  assign Mem1_ext_R0_en = 1'h1;
  assign Mem1_ext_R0_addr = R0_addr;
  assign R0_data = Mem1_ext_R0_data;
  assign Mem1_ext_W0_clk = W0_clk;
  assign Mem1_ext_W0_en = W0_en;
  assign Mem1_ext_W0_addr = W0_addr;
  assign Mem1_ext_W0_data = W0_data;
endmodule
module Mem2(
  input  [7:0]   R0_addr,
  input          R0_clk,
  output [127:0] R0_data,
  input  [7:0]   W0_addr,
  input          W0_en,
  input          W0_clk,
  input  [127:0] W0_data
);
  wire [7:0] Mem2_ext_R0_addr;
  wire  Mem2_ext_R0_en;
  wire  Mem2_ext_R0_clk;
  wire [127:0] Mem2_ext_R0_data;
  wire [7:0] Mem2_ext_W0_addr;
  wire  Mem2_ext_W0_en;
  wire  Mem2_ext_W0_clk;
  wire [127:0] Mem2_ext_W0_data;
  Mem2_ext Mem2_ext (
    .R0_addr(Mem2_ext_R0_addr),
    .R0_en(Mem2_ext_R0_en),
    .R0_clk(Mem2_ext_R0_clk),
    .R0_data(Mem2_ext_R0_data),
    .W0_addr(Mem2_ext_W0_addr),
    .W0_en(Mem2_ext_W0_en),
    .W0_clk(Mem2_ext_W0_clk),
    .W0_data(Mem2_ext_W0_data)
  );
  assign Mem2_ext_R0_clk = R0_clk;
  assign Mem2_ext_R0_en = 1'h1;
  assign Mem2_ext_R0_addr = R0_addr;
  assign R0_data = Mem2_ext_R0_data;
  assign Mem2_ext_W0_clk = W0_clk;
  assign Mem2_ext_W0_en = W0_en;
  assign Mem2_ext_W0_addr = W0_addr;
  assign Mem2_ext_W0_data = W0_data;
endmodule
